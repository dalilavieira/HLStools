-- ----------------------------------------------------------------------------
-- LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
-- Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
-- For technical issues, please contact: support@legupcomputing.com
-- For general inquiries, please contact: info@legupcomputing.com
-- Date: Wed Apr 29 09:18:45 2020
-- ----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

-- LegUp generic types
package legup_types_pkg is
type slv_array_t is array (natural range <> ) of std_logic_vector;

end package legup_types_pkg;

package body legup_types_pkg is
end package body legup_types_pkg;
