library verilog;
use verilog.vl_types.all;
entity legup_pthreadcall_mandelbrot is
    generic(
        LEGUP_0         : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_1: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_2: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_3: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi1);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_4: vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb5_preheader_lr_ph_i_5: vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi1);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb1_i_6: vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi0);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb1_i_7: vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi1);
        LEGUP_loop_pipeline_wait_loop_2_8: vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi0);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb4_i_9: vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi1);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb4_i_10: vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi1, Hi0);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb6_i_11: vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi1, Hi1);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb5_preheader_i_12: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi0, Hi0);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb7_bb8_crit_edge_i_13: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi0, Hi1);
        LEGUP_F_legup_pthreadcall_mandelbrot_BB_mandelbrot_exit_14: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi0)
    );
    port(
        clk             : in     vl_logic;
        clk2x           : in     vl_logic;
        clk1x_follower  : in     vl_logic;
        reset           : in     vl_logic;
        start           : in     vl_logic;
        finish          : out    vl_logic;
        memory_controller_enable_a: out    vl_logic;
        memory_controller_address_a: out    vl_logic_vector(31 downto 0);
        memory_controller_write_enable_a: out    vl_logic;
        memory_controller_in_a: out    vl_logic_vector(63 downto 0);
        memory_controller_size_a: out    vl_logic_vector(1 downto 0);
        memory_controller_out_a: in     vl_logic_vector(63 downto 0);
        memory_controller_enable_b: out    vl_logic;
        memory_controller_address_b: out    vl_logic_vector(31 downto 0);
        memory_controller_write_enable_b: out    vl_logic;
        memory_controller_in_b: out    vl_logic_vector(63 downto 0);
        memory_controller_size_b: out    vl_logic_vector(1 downto 0);
        memory_controller_out_b: in     vl_logic_vector(63 downto 0);
        memory_controller_waitrequest: in     vl_logic;
        return_val      : out    vl_logic_vector(31 downto 0);
        arg_threadarg   : in     vl_logic_vector(31 downto 0);
        arg_threadID    : in     vl_logic_vector(31 downto 0);
        arg_threadIDValue: in     vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LEGUP_0 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_1 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_2 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_3 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_0_4 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb5_preheader_lr_ph_i_5 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb1_i_6 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb1_i_7 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_loop_pipeline_wait_loop_2_8 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb4_i_9 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb4_i_10 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb6_i_11 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb5_preheader_i_12 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_bb7_bb8_crit_edge_i_13 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_legup_pthreadcall_mandelbrot_BB_mandelbrot_exit_14 : constant is 2;
end legup_pthreadcall_mandelbrot;
