// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Mon May  4 13:23:04 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [3:0] LEGUP_0 = 4'd0;
parameter [3:0] LEGUP_F_main_BB_entry_1 = 4'd1;
parameter [3:0] LEGUP_F_main_BB_for_body_2 = 4'd2;
parameter [3:0] LEGUP_F_main_BB_for_body_3 = 4'd3;
parameter [3:0] LEGUP_F_main_BB_for_body_i_preheader_4 = 4'd4;
parameter [3:0] LEGUP_F_main_BB_for_body_i_5 = 4'd5;
parameter [3:0] LEGUP_F_main_BB_for_body_i_6 = 4'd6;
parameter [3:0] LEGUP_F_main_BB_for_body_i_7 = 4'd7;
parameter [3:0] LEGUP_F_main_BB_for_body8_preheader_8 = 4'd8;
parameter [3:0] LEGUP_F_main_BB_for_body8_9 = 4'd9;
parameter [3:0] LEGUP_F_main_BB_for_body8_10 = 4'd10;
parameter [3:0] LEGUP_F_main_BB_for_end14_11 = 4'd11;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [3:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [3:0] next_state;
wire  fsm_stall;
reg [6:0] main_for_body_0;
reg [6:0] main_for_body_0_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_arrayidx;
reg [8:0] main_for_body_sub;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_arrayidx3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_arrayidx4;
reg [7:0] main_for_body_1;
reg [7:0] main_for_body_1_reg;
reg  main_for_body_exitcond2;
reg  main_for_body_exitcond2_reg;
reg [6:0] main_for_body_i_i_08_i;
reg [6:0] main_for_body_i_i_08_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx1_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx2_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx2_i_reg;
reg [31:0] main_for_body_i_2;
reg [31:0] main_for_body_i_3;
reg [31:0] main_for_body_i_add_i;
reg [7:0] main_for_body_i_4;
reg [7:0] main_for_body_i_4_reg;
reg  main_for_body_i_exitcond1;
reg  main_for_body_i_exitcond1_reg;
reg [6:0] main_for_body8_i5_034;
reg [6:0] main_for_body8_i5_034_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body8_arrayidx9;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body8_arrayidx10;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body8_arrayidx11;
reg [31:0] main_for_body8_5;
reg [31:0] main_for_body8_6;
reg [31:0] main_for_body8_7;
reg [7:0] main_for_body8_8;
reg [7:0] main_for_body8_8_reg;
reg  main_for_body8_exitcond;
reg  main_for_body8_exitcond_reg;
reg [6:0] main_entry_vla31_address_a;
reg  main_entry_vla31_write_enable_a;
reg [31:0] main_entry_vla31_in_a;
wire [31:0] main_entry_vla31_out_a;
reg [6:0] main_entry_vla132_address_a;
reg  main_entry_vla132_write_enable_a;
reg [31:0] main_entry_vla132_in_a;
wire [31:0] main_entry_vla132_out_a;
reg [6:0] main_entry_vla233_address_a;
reg  main_entry_vla233_write_enable_a;
reg [31:0] main_entry_vla233_in_a;
wire [31:0] main_entry_vla233_out_a;



//   %vla31 = alloca [100 x i32], align 4, !dbg !35, !MSB !36, !LSB !37, !extendFrom !36
ram_single_port_intel main_entry_vla31 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla31_address_a ),
	.wren_a( main_entry_vla31_write_enable_a ),
	.data_a( main_entry_vla31_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla31_out_a )
);
defparam main_entry_vla31.width_a = 32;
defparam main_entry_vla31.widthad_a = 7;
defparam main_entry_vla31.width_be_a = 4;
defparam main_entry_vla31.numwords_a = 100;
defparam main_entry_vla31.latency = 1;


//   %vla132 = alloca [100 x i32], align 4, !dbg !35, !MSB !36, !LSB !37, !extendFrom !36
ram_single_port_intel main_entry_vla132 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla132_address_a ),
	.wren_a( main_entry_vla132_write_enable_a ),
	.data_a( main_entry_vla132_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla132_out_a )
);
defparam main_entry_vla132.width_a = 32;
defparam main_entry_vla132.widthad_a = 7;
defparam main_entry_vla132.width_be_a = 4;
defparam main_entry_vla132.numwords_a = 100;
defparam main_entry_vla132.latency = 1;


//   %vla233 = alloca [100 x i32], align 4, !dbg !35, !MSB !36, !LSB !37, !extendFrom !36
ram_single_port_intel main_entry_vla233 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla233_address_a ),
	.wren_a( main_entry_vla233_write_enable_a ),
	.data_a( main_entry_vla233_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla233_out_a )
);
defparam main_entry_vla233.width_a = 32;
defparam main_entry_vla233.widthad_a = 7;
defparam main_entry_vla233.width_be_a = 4;
defparam main_entry_vla233.numwords_a = 100;
defparam main_entry_vla233.latency = 1;

/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_for_body8_10)) begin
		$write("%d + %d = %d\n", $signed(main_for_body8_5), $signed(main_for_body8_6), $signed(main_for_body8_7));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_for_body8_5) === 1'bX) finish <= 0;
		if (reset == 1'b0 && ^(main_for_body8_6) === 1'bX) finish <= 0;
		if (reset == 1'b0 && ^(main_for_body8_7) === 1'bX) finish <= 0;
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_for_body_2;
LEGUP_F_main_BB_for_body8_10:
	if ((fsm_stall == 1'd0) && (main_for_body8_exitcond_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_end14_11;
	else if ((fsm_stall == 1'd0) && (main_for_body8_exitcond_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body8_9;
LEGUP_F_main_BB_for_body8_9:
		next_state = LEGUP_F_main_BB_for_body8_10;
LEGUP_F_main_BB_for_body8_preheader_8:
		next_state = LEGUP_F_main_BB_for_body8_9;
LEGUP_F_main_BB_for_body_2:
		next_state = LEGUP_F_main_BB_for_body_3;
LEGUP_F_main_BB_for_body_3:
	if ((fsm_stall == 1'd0) && (main_for_body_exitcond2_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_body_i_preheader_4;
	else if ((fsm_stall == 1'd0) && (main_for_body_exitcond2_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_2;
LEGUP_F_main_BB_for_body_i_5:
		next_state = LEGUP_F_main_BB_for_body_i_6;
LEGUP_F_main_BB_for_body_i_6:
		next_state = LEGUP_F_main_BB_for_body_i_7;
LEGUP_F_main_BB_for_body_i_7:
	if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond1_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_body8_preheader_8;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond1_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_5;
LEGUP_F_main_BB_for_body_i_preheader_4:
		next_state = LEGUP_F_main_BB_for_body_i_5;
LEGUP_F_main_BB_for_end14_11:
		next_state = LEGUP_0;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_0 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_3) & (fsm_stall == 1'd0)) & (main_for_body_exitcond2_reg == 1'd0))) */ begin
		main_for_body_0 = main_for_body_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_0_reg <= main_for_body_0;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_3) & (fsm_stall == 1'd0)) & (main_for_body_exitcond2_reg == 1'd0))) begin
		main_for_body_0_reg <= main_for_body_0;
	end
end
always @(*) begin
		main_for_body_arrayidx = (1'd0 + (4 * {25'd0,main_for_body_0_reg}));
end
always @(*) begin
		main_for_body_sub = (32'd100 - {2'd0,main_for_body_0_reg});
end
always @(*) begin
		main_for_body_arrayidx3 = (1'd0 + (4 * {25'd0,main_for_body_0_reg}));
end
always @(*) begin
		main_for_body_arrayidx4 = (1'd0 + (4 * {25'd0,main_for_body_0_reg}));
end
always @(*) begin
		main_for_body_1 = ({1'd0,main_for_body_0_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_for_body_1_reg <= main_for_body_1;
	end
end
always @(*) begin
		main_for_body_exitcond2 = (main_for_body_1 == 32'd100);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_for_body_exitcond2_reg <= main_for_body_exitcond2;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_08_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_i_7) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond1_reg == 1'd0))) */ begin
		main_for_body_i_i_08_i = main_for_body_i_4_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_08_i_reg <= main_for_body_i_i_08_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_7) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond1_reg == 1'd0))) begin
		main_for_body_i_i_08_i_reg <= main_for_body_i_i_08_i;
	end
end
always @(*) begin
		main_for_body_i_arrayidx_i = (1'd0 + (4 * {25'd0,main_for_body_i_i_08_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx1_i = (1'd0 + (4 * {25'd0,main_for_body_i_i_08_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx2_i = (1'd0 + (4 * {25'd0,main_for_body_i_i_08_i_reg}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_5)) begin
		main_for_body_i_arrayidx2_i_reg <= main_for_body_i_arrayidx2_i;
	end
end
always @(*) begin
		main_for_body_i_2 = main_entry_vla31_out_a;
end
always @(*) begin
		main_for_body_i_3 = main_entry_vla132_out_a;
end
always @(*) begin
		main_for_body_i_add_i = (main_for_body_i_3 + main_for_body_i_2);
end
always @(*) begin
		main_for_body_i_4 = ({1'd0,main_for_body_i_i_08_i_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_5)) begin
		main_for_body_i_4_reg <= main_for_body_i_4;
	end
end
always @(*) begin
		main_for_body_i_exitcond1 = (main_for_body_i_4 == 32'd100);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_5)) begin
		main_for_body_i_exitcond1_reg <= main_for_body_i_exitcond1;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body8_preheader_8) & (fsm_stall == 1'd0))) begin
		main_for_body8_i5_034 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body8_10) & (fsm_stall == 1'd0)) & (main_for_body8_exitcond_reg == 1'd0))) */ begin
		main_for_body8_i5_034 = main_for_body8_8_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body8_preheader_8) & (fsm_stall == 1'd0))) begin
		main_for_body8_i5_034_reg <= main_for_body8_i5_034;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body8_10) & (fsm_stall == 1'd0)) & (main_for_body8_exitcond_reg == 1'd0))) begin
		main_for_body8_i5_034_reg <= main_for_body8_i5_034;
	end
end
always @(*) begin
		main_for_body8_arrayidx9 = (1'd0 + (4 * {25'd0,main_for_body8_i5_034_reg}));
end
always @(*) begin
		main_for_body8_arrayidx10 = (1'd0 + (4 * {25'd0,main_for_body8_i5_034_reg}));
end
always @(*) begin
		main_for_body8_arrayidx11 = (1'd0 + (4 * {25'd0,main_for_body8_i5_034_reg}));
end
always @(*) begin
		main_for_body8_5 = main_entry_vla31_out_a;
end
always @(*) begin
		main_for_body8_6 = main_entry_vla132_out_a;
end
always @(*) begin
		main_for_body8_7 = main_entry_vla233_out_a;
end
always @(*) begin
		main_for_body8_8 = ({1'd0,main_for_body8_i5_034_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body8_9)) begin
		main_for_body8_8_reg <= main_for_body8_8;
	end
end
always @(*) begin
		main_for_body8_exitcond = (main_for_body8_8 == 32'd100);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body8_9)) begin
		main_for_body8_exitcond_reg <= main_for_body8_exitcond;
	end
end
always @(*) begin
	main_entry_vla31_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla31_address_a = (main_for_body_arrayidx >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_5)) begin
		main_entry_vla31_address_a = (main_for_body_i_arrayidx_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body8_9)) begin
		main_entry_vla31_address_a = (main_for_body8_arrayidx9 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla31_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla31_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla31_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla31_in_a = {25'd0,main_for_body_0_reg};
	end
end
always @(*) begin
	main_entry_vla132_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla132_address_a = (main_for_body_arrayidx3 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_5)) begin
		main_entry_vla132_address_a = (main_for_body_i_arrayidx1_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body8_9)) begin
		main_entry_vla132_address_a = (main_for_body8_arrayidx10 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla132_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla132_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla132_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla132_in_a = {{23{main_for_body_sub[8]}},main_for_body_sub};
	end
end
always @(*) begin
	main_entry_vla233_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla233_address_a = (main_for_body_arrayidx4 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_6)) begin
		main_entry_vla233_address_a = (main_for_body_i_arrayidx2_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body8_9)) begin
		main_entry_vla233_address_a = (main_for_body8_arrayidx11 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla233_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla233_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_6)) begin
		main_entry_vla233_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla233_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_vla233_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_6)) begin
		main_entry_vla233_in_a = main_for_body_i_add_i;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end14_11)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end14_11)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
