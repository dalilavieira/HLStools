library verilog;
use verilog.vl_types.all;
entity fadd64_altbarrel_shift_95g is
    port(
        aclr            : in     vl_logic;
        clk_en          : in     vl_logic;
        clock           : in     vl_logic;
        data            : in     vl_logic_vector(54 downto 0);
        distance        : in     vl_logic_vector(5 downto 0);
        result          : out    vl_logic_vector(54 downto 0)
    );
end fadd64_altbarrel_shift_95g;
