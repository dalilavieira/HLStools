// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Mon Apr 20 08:57:44 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [3:0] LEGUP_0 = 4'd0;
parameter [3:0] LEGUP_F_main_BB_entry_1 = 4'd1;
parameter [3:0] LEGUP_F_main_BB_for_body_i_2 = 4'd2;
parameter [3:0] LEGUP_F_main_BB_for_body_i_3 = 4'd3;
parameter [3:0] LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4 = 4'd4;
parameter [3:0] LEGUP_F_main_BB_for_cond10_preheader_i_5 = 4'd5;
parameter [3:0] LEGUP_F_main_BB_for_body13_i_6 = 4'd6;
parameter [3:0] LEGUP_F_main_BB_for_body13_i_7 = 4'd7;
parameter [3:0] LEGUP_F_main_BB_for_body13_i_8 = 4'd8;
parameter [3:0] LEGUP_F_main_BB_for_body13_i_9 = 4'd9;
parameter [3:0] LEGUP_F_main_BB_for_body13_i_10 = 4'd10;
parameter [3:0] LEGUP_F_main_BB_for_body13_i_11 = 4'd11;
parameter [3:0] LEGUP_F_main_BB_for_body13_i_12 = 4'd12;
parameter [3:0] LEGUP_F_main_BB_for_inc113_i_13 = 4'd13;
parameter [3:0] LEGUP_F_main_BB_poly6_exit_14 = 4'd14;
parameter [3:0] LEGUP_F_main_BB_poly6_exit_15 = 4'd15;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [3:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [3:0] next_state;
wire  fsm_stall;
reg [10:0] main_for_body_i_k_0162_i;
reg [10:0] main_for_body_i_k_0162_i_reg;
reg [15:0] main_for_body_i_bit_select17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx2_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx4_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx5_i;
reg [11:0] main_for_body_i_0;
reg [11:0] main_for_body_i_0_reg;
reg  main_for_body_i_exitcond5;
reg  main_for_body_i_exitcond5_reg;
reg [6:0] main_for_cond10_preheader_i_i_0161_i;
reg [6:0] main_for_cond10_preheader_i_i_0161_i_reg;
reg [31:0] main_for_body13_i_k_1160_i;
reg [31:0] main_for_body13_i_k_1160_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx14_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx16_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx30_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx109_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx109_i_reg;
reg [15:0] main_for_body13_i_1;
reg [31:0] main_for_body13_i_bit_concat16;
reg [15:0] main_for_body13_i_2;
reg [31:0] main_for_body13_i_bit_concat15;
reg [31:0] main_for_body13_i_bit_concat15_reg;
reg [31:0] main_for_body13_i_bit_concat14;
reg [31:0] main_for_body13_i_tmp_i;
reg [31:0] main_for_body13_i_mul25_i;
reg [15:0] main_for_body13_i_3;
reg [31:0] main_for_body13_i_bit_concat13;
reg [31:0] main_for_body13_i_bit_concat13_reg;
reg [31:0] main_for_body13_i_mul36_i;
reg [31:0] main_for_body13_i_mul39_i;
reg [31:0] main_for_body13_i_bit_concat12;
reg [31:0] main_for_body13_i_bit_concat11;
reg [31:0] main_for_body13_i_sr_add7;
reg [31:0] main_for_body13_i_sub_i;
reg [31:0] main_for_body13_i_sub_i_reg;
reg [31:0] main_for_body13_i_mul47_i;
reg [31:0] main_for_body13_i_sr_negate;
reg [30:0] main_for_body13_i_bit_select9;
reg [31:0] main_for_body13_i_bit_concat10;
reg [31:0] main_for_body13_i_bit_concat8;
reg [31:0] main_for_body13_i_sr_add8;
reg [31:0] main_for_body13_i_bit_concat7;
reg [31:0] main_for_body13_i_bit_concat6;
reg [31:0] main_for_body13_i_sr_add10;
reg [31:0] main_for_body13_i_sr_add10_reg;
reg [31:0] main_for_body13_i_newEarly_sub53_i;
reg [31:0] main_for_body13_i_newEarly_sub53_i_reg;
reg [31:0] main_for_body13_i_newCurOp_sub53_i;
reg [31:0] main_for_body13_i_mul54_i;
reg [31:0] main_for_body13_i_mul54_i_reg;
reg [31:0] main_for_body13_i_sub55_i;
reg [31:0] main_for_body13_i_bit_concat5;
reg [31:0] main_for_body13_i_bit_concat4;
reg [31:0] main_for_body13_i_sr_add13;
reg [31:0] main_for_body13_i_newEarly_sub61_i;
reg [31:0] main_for_body13_i_newCurOp_sub61_i;
reg [31:0] main_for_body13_i_mul62_i;
reg [31:0] main_for_body13_i_mul62_i_reg;
reg [31:0] main_for_body13_i_sub63_i;
reg [31:0] main_for_body13_i_sub75_i;
reg [31:0] main_for_body13_i_mul76_i;
reg [31:0] main_for_body13_i_sub81_i;
reg [31:0] main_for_body13_i_mul82_i;
reg [31:0] main_for_body13_i_add83_i;
reg [31:0] main_for_body13_i_mul84_i;
reg [31:0] main_for_body13_i_sr_negate14;
reg [31:0] main_for_body13_i_bit_concat3;
reg [31:0] main_for_body13_i_sr_add17;
reg [31:0] main_for_body13_i_bit_concat2;
reg [31:0] main_for_body13_i_bit_concat1;
reg [31:0] main_for_body13_i_sr_add20;
reg [31:0] main_for_body13_i_sr_add20_reg;
reg [31:0] main_for_body13_i_newEarly_add90_i;
reg [31:0] main_for_body13_i_newEarly_add90_i_reg;
reg [31:0] main_for_body13_i_newCurOp_add90_i;
reg [31:0] main_for_body13_i_mul91_i;
reg [31:0] main_for_body13_i_sub92_i;
reg [31:0] main_for_body13_i_sub99_i;
reg [31:0] main_for_body13_i_mul100_i;
reg [31:0] main_for_body13_i_sub101_i;
reg [31:0] main_for_body13_i_mul102_i;
reg [31:0] main_for_body13_i_add103_i;
reg [31:0] main_for_body13_i_mul104_i;
reg [31:0] main_for_body13_i_sub105_i;
reg [31:0] main_for_body13_i_mul106_i;
reg [31:0] main_for_body13_i_tmp158_i;
reg [31:0] main_for_body13_i_tmp159_i;
reg [31:0] main_for_body13_i_tmp159_i_reg;
reg [31:0] main_for_body13_i_sub107_i;
reg [15:0] main_for_body13_i_bit_select;
reg [31:0] main_for_body13_i_4;
reg [31:0] main_for_body13_i_4_reg;
reg  main_for_body13_i_exitcond3;
reg  main_for_body13_i_exitcond3_reg;
reg [7:0] main_for_inc113_i_5;
reg  main_for_inc113_i_exitcond4;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_poly6_exit_arrayidx116_i;
reg [15:0] main_poly6_exit_6;
reg [31:0] main_poly6_exit_bit_concat;
reg [9:0] main_entry_a_i_address_a;
reg  main_entry_a_i_write_enable_a;
reg [15:0] main_entry_a_i_in_a;
wire [15:0] main_entry_a_i_out_a;
reg [9:0] main_entry_b_i_address_a;
reg  main_entry_b_i_write_enable_a;
reg [15:0] main_entry_b_i_in_a;
wire [15:0] main_entry_b_i_out_a;
reg [9:0] main_entry_c_i_address_a;
reg  main_entry_c_i_write_enable_a;
reg [15:0] main_entry_c_i_in_a;
wire [15:0] main_entry_c_i_out_a;
reg [9:0] main_entry_out_i_address_a;
reg  main_entry_out_i_write_enable_a;
reg [15:0] main_entry_out_i_in_a;
wire [15:0] main_entry_out_i_out_a;
reg [15:0] main_for_body_i_k_0162_i_reg_width_extended;
wire [15:0] main_for_body13_i_bit_concat16_bit_select_operand_0;
wire [15:0] main_for_body13_i_bit_concat15_bit_select_operand_0;
wire [12:0] main_for_body13_i_bit_concat14_bit_select_operand_0;
wire [2:0] main_for_body13_i_bit_concat14_bit_select_operand_4;
reg  legup_mult_main_for_body13_i_mul25_i_en;
reg [31:0] main_for_body13_i_mul25_i_stage0_reg;
wire [15:0] main_for_body13_i_bit_concat13_bit_select_operand_0;
reg  legup_mult_main_for_body13_i_mul36_i_en;
reg [31:0] main_for_body13_i_mul36_i_stage0_reg;
wire [14:0] main_for_body13_i_bit_concat12_bit_select_operand_0;
wire  main_for_body13_i_bit_concat12_bit_select_operand_4;
wire [12:0] main_for_body13_i_bit_concat11_bit_select_operand_0;
wire [2:0] main_for_body13_i_bit_concat11_bit_select_operand_4;
wire  main_for_body13_i_bit_concat10_bit_select_operand_2;
wire [10:0] main_for_body13_i_bit_concat8_bit_select_operand_0;
wire [4:0] main_for_body13_i_bit_concat8_bit_select_operand_4;
wire [8:0] main_for_body13_i_bit_concat7_bit_select_operand_0;
wire [6:0] main_for_body13_i_bit_concat7_bit_select_operand_4;
wire [7:0] main_for_body13_i_bit_concat6_bit_select_operand_0;
wire [7:0] main_for_body13_i_bit_concat6_bit_select_operand_4;
wire [5:0] main_for_body13_i_bit_concat5_bit_select_operand_0;
wire [9:0] main_for_body13_i_bit_concat5_bit_select_operand_4;
wire [4:0] main_for_body13_i_bit_concat4_bit_select_operand_0;
wire [10:0] main_for_body13_i_bit_concat4_bit_select_operand_4;
reg  legup_mult_main_for_body13_i_mul62_i_en;
reg [31:0] main_for_body13_i_mul62_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul76_i_en;
reg [31:0] main_for_body13_i_mul76_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul82_i_en;
reg [31:0] main_for_body13_i_mul82_i_stage0_reg;
wire [12:0] main_for_body13_i_bit_concat3_bit_select_operand_0;
wire [2:0] main_for_body13_i_bit_concat3_bit_select_operand_4;
wire [11:0] main_for_body13_i_bit_concat2_bit_select_operand_0;
wire [3:0] main_for_body13_i_bit_concat2_bit_select_operand_4;
wire [9:0] main_for_body13_i_bit_concat1_bit_select_operand_0;
wire [5:0] main_for_body13_i_bit_concat1_bit_select_operand_4;
reg  legup_mult_main_for_body13_i_mul100_i_en;
reg [31:0] main_for_body13_i_mul100_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul39_i_en;
reg [31:0] main_for_body13_i_mul39_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul54_i_en;
reg [31:0] main_for_body13_i_mul54_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul84_i_en;
reg [31:0] main_for_body13_i_mul84_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul91_i_en;
reg [31:0] main_for_body13_i_mul91_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul102_i_en;
reg [31:0] main_for_body13_i_mul102_i_stage0_reg;
reg  legup_mult_main_for_body13_i_tmp159_i_en;
reg [31:0] main_for_body13_i_tmp159_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul47_i_en;
reg [31:0] main_for_body13_i_mul47_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul104_i_en;
reg [31:0] main_for_body13_i_mul104_i_stage0_reg;
reg  legup_mult_main_for_body13_i_mul106_i_en;
reg [31:0] main_for_body13_i_mul106_i_stage0_reg;
wire [15:0] main_poly6_exit_bit_concat_bit_select_operand_0;



//   %a.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port_intel main_entry_a_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_a_i_address_a ),
	.wren_a( main_entry_a_i_write_enable_a ),
	.data_a( main_entry_a_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_a_i_out_a )
);
defparam main_entry_a_i.width_a = 16;
defparam main_entry_a_i.widthad_a = 10;
defparam main_entry_a_i.width_be_a = 2;
defparam main_entry_a_i.numwords_a = 1024;
defparam main_entry_a_i.latency = 1;


//   %b.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port_intel main_entry_b_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_b_i_address_a ),
	.wren_a( main_entry_b_i_write_enable_a ),
	.data_a( main_entry_b_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_b_i_out_a )
);
defparam main_entry_b_i.width_a = 16;
defparam main_entry_b_i.widthad_a = 10;
defparam main_entry_b_i.width_be_a = 2;
defparam main_entry_b_i.numwords_a = 1024;
defparam main_entry_b_i.latency = 1;


//   %c.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port_intel main_entry_c_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_c_i_address_a ),
	.wren_a( main_entry_c_i_write_enable_a ),
	.data_a( main_entry_c_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_c_i_out_a )
);
defparam main_entry_c_i.width_a = 16;
defparam main_entry_c_i.widthad_a = 10;
defparam main_entry_c_i.width_be_a = 2;
defparam main_entry_c_i.numwords_a = 1024;
defparam main_entry_c_i.latency = 1;


//   %out.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port_intel main_entry_out_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_out_i_address_a ),
	.wren_a( main_entry_out_i_write_enable_a ),
	.data_a( main_entry_out_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_out_i_out_a )
);
defparam main_entry_out_i.width_a = 16;
defparam main_entry_out_i.widthad_a = 10;
defparam main_entry_out_i.width_be_a = 2;
defparam main_entry_out_i.numwords_a = 1024;
defparam main_entry_out_i.latency = 1;

/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_poly6_exit_15)) begin
		$write("%d\n", $signed(main_poly6_exit_bit_concat));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_poly6_exit_bit_concat) === 1'bX) finish <= 0;
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_for_body_i_2;
LEGUP_F_main_BB_for_body13_i_10:
		next_state = LEGUP_F_main_BB_for_body13_i_11;
LEGUP_F_main_BB_for_body13_i_11:
		next_state = LEGUP_F_main_BB_for_body13_i_12;
LEGUP_F_main_BB_for_body13_i_12:
	if ((fsm_stall == 1'd0) && (main_for_body13_i_exitcond3_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc113_i_13;
	else if ((fsm_stall == 1'd0) && (main_for_body13_i_exitcond3_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body13_i_6;
LEGUP_F_main_BB_for_body13_i_6:
		next_state = LEGUP_F_main_BB_for_body13_i_7;
LEGUP_F_main_BB_for_body13_i_7:
		next_state = LEGUP_F_main_BB_for_body13_i_8;
LEGUP_F_main_BB_for_body13_i_8:
		next_state = LEGUP_F_main_BB_for_body13_i_9;
LEGUP_F_main_BB_for_body13_i_9:
		next_state = LEGUP_F_main_BB_for_body13_i_10;
LEGUP_F_main_BB_for_body_i_2:
		next_state = LEGUP_F_main_BB_for_body_i_3;
LEGUP_F_main_BB_for_body_i_3:
	if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond5_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond5_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_2;
LEGUP_F_main_BB_for_cond10_preheader_i_5:
		next_state = LEGUP_F_main_BB_for_body13_i_6;
LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4:
		next_state = LEGUP_F_main_BB_for_cond10_preheader_i_5;
LEGUP_F_main_BB_for_inc113_i_13:
	if ((fsm_stall == 1'd0) && (main_for_inc113_i_exitcond4 == 1'd1))
		next_state = LEGUP_F_main_BB_poly6_exit_14;
	else if ((fsm_stall == 1'd0) && (main_for_inc113_i_exitcond4 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond10_preheader_i_5;
LEGUP_F_main_BB_poly6_exit_14:
		next_state = LEGUP_F_main_BB_poly6_exit_15;
LEGUP_F_main_BB_poly6_exit_15:
		next_state = LEGUP_0;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_i_k_0162_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_i_3) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond5_reg == 1'd0))) */ begin
		main_for_body_i_k_0162_i = main_for_body_i_0_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_i_k_0162_i_reg <= main_for_body_i_k_0162_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_3) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond5_reg == 1'd0))) begin
		main_for_body_i_k_0162_i_reg <= main_for_body_i_k_0162_i;
	end
end
always @(*) begin
		main_for_body_i_bit_select17 = main_for_body_i_k_0162_i_reg_width_extended[15:0];
end
always @(*) begin
		main_for_body_i_arrayidx_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0162_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx2_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0162_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx4_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0162_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx5_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0162_i_reg}));
end
always @(*) begin
		main_for_body_i_0 = ({1'd0,main_for_body_i_k_0162_i_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_for_body_i_0_reg <= main_for_body_i_0;
	end
end
always @(*) begin
		main_for_body_i_exitcond5 = (main_for_body_i_0 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_for_body_i_exitcond5_reg <= main_for_body_i_exitcond5;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_cond10_preheader_i_i_0161_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc113_i_13) & (fsm_stall == 1'd0)) & (main_for_inc113_i_exitcond4 == 1'd0))) */ begin
		main_for_cond10_preheader_i_i_0161_i = main_for_inc113_i_5;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_cond10_preheader_i_i_0161_i_reg <= main_for_cond10_preheader_i_i_0161_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc113_i_13) & (fsm_stall == 1'd0)) & (main_for_inc113_i_exitcond4 == 1'd0))) begin
		main_for_cond10_preheader_i_i_0161_i_reg <= main_for_cond10_preheader_i_i_0161_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_5) & (fsm_stall == 1'd0))) begin
		main_for_body13_i_k_1160_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body13_i_12) & (fsm_stall == 1'd0)) & (main_for_body13_i_exitcond3_reg == 1'd0))) */ begin
		main_for_body13_i_k_1160_i = main_for_body13_i_4_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_5) & (fsm_stall == 1'd0))) begin
		main_for_body13_i_k_1160_i_reg <= main_for_body13_i_k_1160_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body13_i_12) & (fsm_stall == 1'd0)) & (main_for_body13_i_exitcond3_reg == 1'd0))) begin
		main_for_body13_i_k_1160_i_reg <= main_for_body13_i_k_1160_i;
	end
end
always @(*) begin
		main_for_body13_i_arrayidx14_i = (1'd0 + (2 * main_for_body13_i_k_1160_i_reg));
end
always @(*) begin
		main_for_body13_i_arrayidx16_i = (1'd0 + (2 * main_for_body13_i_k_1160_i_reg));
end
always @(*) begin
		main_for_body13_i_arrayidx30_i = (1'd0 + (2 * main_for_body13_i_k_1160_i_reg));
end
always @(*) begin
		main_for_body13_i_arrayidx109_i = (1'd0 + (2 * main_for_body13_i_k_1160_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_for_body13_i_arrayidx109_i_reg <= main_for_body13_i_arrayidx109_i;
	end
end
always @(*) begin
		main_for_body13_i_1 = main_entry_b_i_out_a;
end
always @(*) begin
		main_for_body13_i_bit_concat16 = {main_for_body13_i_bit_concat16_bit_select_operand_0[15:0], main_for_body13_i_1[15:0]};
end
always @(*) begin
		main_for_body13_i_2 = main_entry_c_i_out_a;
end
always @(*) begin
		main_for_body13_i_bit_concat15 = {main_for_body13_i_bit_concat15_bit_select_operand_0[15:0], main_for_body13_i_2[15:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_bit_concat15_reg <= main_for_body13_i_bit_concat15;
	end
end
always @(*) begin
		main_for_body13_i_bit_concat14 = {{main_for_body13_i_bit_concat14_bit_select_operand_0[12:0], main_for_body13_i_1[15:0]}, main_for_body13_i_bit_concat14_bit_select_operand_4[2:0]};
end
always @(*) begin
		main_for_body13_i_tmp_i = (main_for_body13_i_bit_concat14 + 32'd126144);
end
always @(*) begin
	main_for_body13_i_mul25_i = main_for_body13_i_mul25_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_3 = main_entry_a_i_out_a;
end
always @(*) begin
		main_for_body13_i_bit_concat13 = {main_for_body13_i_bit_concat13_bit_select_operand_0[15:0], main_for_body13_i_3[15:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_bit_concat13_reg <= main_for_body13_i_bit_concat13;
	end
end
always @(*) begin
	main_for_body13_i_mul36_i = main_for_body13_i_mul36_i_stage0_reg;
end
always @(*) begin
	main_for_body13_i_mul39_i = main_for_body13_i_mul39_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_bit_concat12 = {{main_for_body13_i_bit_concat12_bit_select_operand_0[14:0], main_for_body13_i_1[15:0]}, main_for_body13_i_bit_concat12_bit_select_operand_4};
end
always @(*) begin
		main_for_body13_i_bit_concat11 = {{main_for_body13_i_bit_concat11_bit_select_operand_0[12:0], main_for_body13_i_1[15:0]}, main_for_body13_i_bit_concat11_bit_select_operand_4[2:0]};
end
always @(*) begin
		main_for_body13_i_sr_add7 = (main_for_body13_i_bit_concat12 + main_for_body13_i_bit_concat11);
end
always @(*) begin
		main_for_body13_i_sub_i = (main_for_body13_i_sr_add7 + $signed(-32'd432));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_sub_i_reg <= main_for_body13_i_sub_i;
	end
end
always @(*) begin
	main_for_body13_i_mul47_i = main_for_body13_i_mul47_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sr_negate = (32'd0 - main_for_body13_i_bit_concat15);
end
always @(*) begin
		main_for_body13_i_bit_select9 = main_for_body13_i_sr_negate[30:0];
end
always @(*) begin
		main_for_body13_i_bit_concat10 = {main_for_body13_i_bit_select9[30:0], main_for_body13_i_bit_concat10_bit_select_operand_2};
end
always @(*) begin
		main_for_body13_i_bit_concat8 = {{main_for_body13_i_bit_concat8_bit_select_operand_0[10:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat8_bit_select_operand_4[4:0]};
end
always @(*) begin
		main_for_body13_i_sr_add8 = (main_for_body13_i_bit_concat10 + main_for_body13_i_bit_concat8);
end
always @(*) begin
		main_for_body13_i_bit_concat7 = {{main_for_body13_i_bit_concat7_bit_select_operand_0[8:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat7_bit_select_operand_4[6:0]};
end
always @(*) begin
		main_for_body13_i_bit_concat6 = {{main_for_body13_i_bit_concat6_bit_select_operand_0[7:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat6_bit_select_operand_4[7:0]};
end
always @(*) begin
		main_for_body13_i_sr_add10 = (main_for_body13_i_bit_concat7 + main_for_body13_i_bit_concat6);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_sr_add10_reg <= main_for_body13_i_sr_add10;
	end
end
always @(*) begin
		main_for_body13_i_newEarly_sub53_i = (main_for_body13_i_sr_add8 + $signed(-32'd20736));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_newEarly_sub53_i_reg <= main_for_body13_i_newEarly_sub53_i;
	end
end
always @(*) begin
		main_for_body13_i_newCurOp_sub53_i = (main_for_body13_i_newEarly_sub53_i_reg + main_for_body13_i_sr_add10_reg);
end
always @(*) begin
	main_for_body13_i_mul54_i = main_for_body13_i_mul54_i_stage0_reg;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_9)) begin
		main_for_body13_i_mul54_i_reg <= main_for_body13_i_mul54_i;
	end
end
always @(*) begin
		main_for_body13_i_sub55_i = (main_for_body13_i_mul47_i - main_for_body13_i_mul54_i_reg);
end
always @(*) begin
		main_for_body13_i_bit_concat5 = {{main_for_body13_i_bit_concat5_bit_select_operand_0[5:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat5_bit_select_operand_4[9:0]};
end
always @(*) begin
		main_for_body13_i_bit_concat4 = {{main_for_body13_i_bit_concat4_bit_select_operand_0[4:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat4_bit_select_operand_4[10:0]};
end
always @(*) begin
		main_for_body13_i_sr_add13 = (main_for_body13_i_bit_concat5 + main_for_body13_i_bit_concat4);
end
always @(*) begin
		main_for_body13_i_newEarly_sub61_i = (main_for_body13_i_sr_add10 + $signed(-32'd1492992));
end
always @(*) begin
		main_for_body13_i_newCurOp_sub61_i = (main_for_body13_i_newEarly_sub61_i + main_for_body13_i_sr_add13);
end
always @(*) begin
	main_for_body13_i_mul62_i = main_for_body13_i_mul62_i_stage0_reg;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_8)) begin
		main_for_body13_i_mul62_i_reg <= main_for_body13_i_mul62_i;
	end
end
always @(*) begin
		main_for_body13_i_sub63_i = (main_for_body13_i_sub55_i - main_for_body13_i_mul62_i_reg);
end
always @(*) begin
		main_for_body13_i_sub75_i = (main_for_body13_i_bit_concat15 + $signed(-32'd32));
end
always @(*) begin
	main_for_body13_i_mul76_i = main_for_body13_i_mul76_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sub81_i = (main_for_body13_i_bit_concat15 + $signed(-32'd72));
end
always @(*) begin
	main_for_body13_i_mul82_i = main_for_body13_i_mul82_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_add83_i = (main_for_body13_i_mul76_i + main_for_body13_i_mul82_i);
end
always @(*) begin
	main_for_body13_i_mul84_i = main_for_body13_i_mul84_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sr_negate14 = (32'd0 - main_for_body13_i_bit_concat15);
end
always @(*) begin
		main_for_body13_i_bit_concat3 = {{main_for_body13_i_bit_concat3_bit_select_operand_0[12:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat3_bit_select_operand_4[2:0]};
end
always @(*) begin
		main_for_body13_i_sr_add17 = (main_for_body13_i_sr_negate14 + main_for_body13_i_bit_concat3);
end
always @(*) begin
		main_for_body13_i_bit_concat2 = {{main_for_body13_i_bit_concat2_bit_select_operand_0[11:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat2_bit_select_operand_4[3:0]};
end
always @(*) begin
		main_for_body13_i_bit_concat1 = {{main_for_body13_i_bit_concat1_bit_select_operand_0[9:0], main_for_body13_i_2[15:0]}, main_for_body13_i_bit_concat1_bit_select_operand_4[5:0]};
end
always @(*) begin
		main_for_body13_i_sr_add20 = (main_for_body13_i_bit_concat2 + main_for_body13_i_bit_concat1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_sr_add20_reg <= main_for_body13_i_sr_add20;
	end
end
always @(*) begin
		main_for_body13_i_newEarly_add90_i = (main_for_body13_i_sr_add17 + 32'd2592);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_newEarly_add90_i_reg <= main_for_body13_i_newEarly_add90_i;
	end
end
always @(*) begin
		main_for_body13_i_newCurOp_add90_i = (main_for_body13_i_newEarly_add90_i_reg + main_for_body13_i_sr_add20_reg);
end
always @(*) begin
	main_for_body13_i_mul91_i = main_for_body13_i_mul91_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sub92_i = (main_for_body13_i_mul84_i - main_for_body13_i_mul91_i);
end
always @(*) begin
		main_for_body13_i_sub99_i = (main_for_body13_i_bit_concat15 + $signed(-32'd864));
end
always @(*) begin
	main_for_body13_i_mul100_i = main_for_body13_i_mul100_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sub101_i = (main_for_body13_i_mul100_i + $signed(-32'd186624));
end
always @(*) begin
	main_for_body13_i_mul102_i = main_for_body13_i_mul102_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_add103_i = (main_for_body13_i_sub92_i + main_for_body13_i_mul102_i);
end
always @(*) begin
	main_for_body13_i_mul104_i = main_for_body13_i_mul104_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sub105_i = (main_for_body13_i_sub63_i - main_for_body13_i_mul104_i);
end
always @(*) begin
	main_for_body13_i_mul106_i = main_for_body13_i_mul106_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_tmp158_i = (main_for_body13_i_mul25_i + 32'd2985984);
end
always @(*) begin
	main_for_body13_i_tmp159_i = main_for_body13_i_tmp159_i_stage0_reg;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_9)) begin
		main_for_body13_i_tmp159_i_reg <= main_for_body13_i_tmp159_i;
	end
end
always @(*) begin
		main_for_body13_i_sub107_i = (main_for_body13_i_tmp159_i_reg - main_for_body13_i_mul106_i);
end
always @(*) begin
		main_for_body13_i_bit_select = main_for_body13_i_sub107_i[15:0];
end
always @(*) begin
		main_for_body13_i_4 = (main_for_body13_i_k_1160_i_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_for_body13_i_4_reg <= main_for_body13_i_4;
	end
end
always @(*) begin
		main_for_body13_i_exitcond3 = (main_for_body13_i_4 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_for_body13_i_exitcond3_reg <= main_for_body13_i_exitcond3;
	end
end
always @(*) begin
		main_for_inc113_i_5 = ({1'd0,main_for_cond10_preheader_i_i_0161_i_reg} + 32'd1);
end
always @(*) begin
		main_for_inc113_i_exitcond4 = (main_for_inc113_i_5 == 32'd100);
end
assign main_poly6_exit_arrayidx116_i = (1'd0 + (2 * 32'd50));
always @(*) begin
		main_poly6_exit_6 = main_entry_out_i_out_a;
end
always @(*) begin
		main_poly6_exit_bit_concat = {main_poly6_exit_bit_concat_bit_select_operand_0[15:0], main_poly6_exit_6[15:0]};
end
always @(*) begin
	main_entry_a_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_a_i_address_a = (main_for_body_i_arrayidx_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_entry_a_i_address_a = (main_for_body13_i_arrayidx30_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_a_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_a_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_a_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_a_i_in_a = main_for_body_i_bit_select17;
	end
end
always @(*) begin
	main_entry_b_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_b_i_address_a = (main_for_body_i_arrayidx2_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_entry_b_i_address_a = (main_for_body13_i_arrayidx14_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_b_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_b_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_b_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_b_i_in_a = main_for_body_i_bit_select17;
	end
end
always @(*) begin
	main_entry_c_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_c_i_address_a = (main_for_body_i_arrayidx4_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_entry_c_i_address_a = (main_for_body13_i_arrayidx16_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_c_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_c_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_c_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_c_i_in_a = main_for_body_i_bit_select17;
	end
end
always @(*) begin
	main_entry_out_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_out_i_address_a = (main_for_body_i_arrayidx5_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_11)) begin
		main_entry_out_i_address_a = (main_for_body13_i_arrayidx109_i_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_poly6_exit_14)) begin
		main_entry_out_i_address_a = (main_poly6_exit_arrayidx116_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_out_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_out_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_11)) begin
		main_entry_out_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_out_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_out_i_in_a = 16'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_11)) begin
		main_entry_out_i_in_a = main_for_body13_i_bit_select;
	end
end
always @(*) begin
	main_for_body_i_k_0162_i_reg_width_extended = {5'd0,main_for_body_i_k_0162_i_reg};
end
assign main_for_body13_i_bit_concat16_bit_select_operand_0 = 16'd0;
assign main_for_body13_i_bit_concat15_bit_select_operand_0 = 16'd0;
assign main_for_body13_i_bit_concat14_bit_select_operand_0 = 13'd0;
assign main_for_body13_i_bit_concat14_bit_select_operand_4 = 3'd0;
always @(*) begin
	legup_mult_main_for_body13_i_mul25_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul25_i_en == 1'd1)) begin
		main_for_body13_i_mul25_i_stage0_reg <= (main_for_body13_i_tmp_i * main_for_body13_i_bit_concat16);
	end
end
assign main_for_body13_i_bit_concat13_bit_select_operand_0 = 16'd0;
always @(*) begin
	legup_mult_main_for_body13_i_mul36_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul36_i_en == 1'd1)) begin
		main_for_body13_i_mul36_i_stage0_reg <= (main_for_body13_i_bit_concat16 * main_for_body13_i_bit_concat16);
	end
end
assign main_for_body13_i_bit_concat12_bit_select_operand_0 = 15'd0;
assign main_for_body13_i_bit_concat12_bit_select_operand_4 = 1'd0;
assign main_for_body13_i_bit_concat11_bit_select_operand_0 = 13'd0;
assign main_for_body13_i_bit_concat11_bit_select_operand_4 = 3'd0;
assign main_for_body13_i_bit_concat10_bit_select_operand_2 = 1'd0;
assign main_for_body13_i_bit_concat8_bit_select_operand_0 = 11'd0;
assign main_for_body13_i_bit_concat8_bit_select_operand_4 = 5'd0;
assign main_for_body13_i_bit_concat7_bit_select_operand_0 = 9'd0;
assign main_for_body13_i_bit_concat7_bit_select_operand_4 = 7'd0;
assign main_for_body13_i_bit_concat6_bit_select_operand_0 = 8'd0;
assign main_for_body13_i_bit_concat6_bit_select_operand_4 = 8'd0;
assign main_for_body13_i_bit_concat5_bit_select_operand_0 = 6'd0;
assign main_for_body13_i_bit_concat5_bit_select_operand_4 = 10'd0;
assign main_for_body13_i_bit_concat4_bit_select_operand_0 = 5'd0;
assign main_for_body13_i_bit_concat4_bit_select_operand_4 = 11'd0;
always @(*) begin
	legup_mult_main_for_body13_i_mul62_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul62_i_en == 1'd1)) begin
		main_for_body13_i_mul62_i_stage0_reg <= (main_for_body13_i_newCurOp_sub61_i * main_for_body13_i_bit_concat15);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul76_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul76_i_en == 1'd1)) begin
		main_for_body13_i_mul76_i_stage0_reg <= (main_for_body13_i_sub75_i * main_for_body13_i_bit_concat16);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul82_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul82_i_en == 1'd1)) begin
		main_for_body13_i_mul82_i_stage0_reg <= (main_for_body13_i_sub81_i * main_for_body13_i_bit_concat15);
	end
end
assign main_for_body13_i_bit_concat3_bit_select_operand_0 = 13'd0;
assign main_for_body13_i_bit_concat3_bit_select_operand_4 = 3'd0;
assign main_for_body13_i_bit_concat2_bit_select_operand_0 = 12'd0;
assign main_for_body13_i_bit_concat2_bit_select_operand_4 = 4'd0;
assign main_for_body13_i_bit_concat1_bit_select_operand_0 = 10'd0;
assign main_for_body13_i_bit_concat1_bit_select_operand_4 = 6'd0;
always @(*) begin
	legup_mult_main_for_body13_i_mul100_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul100_i_en == 1'd1)) begin
		main_for_body13_i_mul100_i_stage0_reg <= (main_for_body13_i_sub99_i * main_for_body13_i_bit_concat15);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul39_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul39_i_en == 1'd1)) begin
		main_for_body13_i_mul39_i_stage0_reg <= (main_for_body13_i_mul36_i * main_for_body13_i_bit_concat15_reg);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul54_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul54_i_en == 1'd1)) begin
		main_for_body13_i_mul54_i_stage0_reg <= (main_for_body13_i_newCurOp_sub53_i * main_for_body13_i_bit_concat15_reg);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul84_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul84_i_en == 1'd1)) begin
		main_for_body13_i_mul84_i_stage0_reg <= (main_for_body13_i_add83_i * main_for_body13_i_mul36_i);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul91_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul91_i_en == 1'd1)) begin
		main_for_body13_i_mul91_i_stage0_reg <= (main_for_body13_i_newCurOp_add90_i * main_for_body13_i_bit_concat15_reg);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul102_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul102_i_en == 1'd1)) begin
		main_for_body13_i_mul102_i_stage0_reg <= (main_for_body13_i_sub101_i * main_for_body13_i_bit_concat15_reg);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_tmp159_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_tmp159_i_en == 1'd1)) begin
		main_for_body13_i_tmp159_i_stage0_reg <= (main_for_body13_i_tmp158_i * main_for_body13_i_bit_concat15_reg);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul47_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul47_i_en == 1'd1)) begin
		main_for_body13_i_mul47_i_stage0_reg <= (main_for_body13_i_mul39_i * main_for_body13_i_sub_i_reg);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul104_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul104_i_en == 1'd1)) begin
		main_for_body13_i_mul104_i_stage0_reg <= (main_for_body13_i_add103_i * main_for_body13_i_bit_concat13_reg);
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul106_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul106_i_en == 1'd1)) begin
		main_for_body13_i_mul106_i_stage0_reg <= (main_for_body13_i_sub105_i * main_for_body13_i_bit_concat13_reg);
	end
end
assign main_poly6_exit_bit_concat_bit_select_operand_0 = 16'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_poly6_exit_15)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_poly6_exit_15)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
