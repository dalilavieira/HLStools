// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Mon Apr 27 08:23:06 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [4:0] LEGUP_0 = 5'd0;
parameter [4:0] LEGUP_F_main_BB_entry_1 = 5'd1;
parameter [4:0] LEGUP_F_main_BB_for_body_i_2 = 5'd2;
parameter [4:0] LEGUP_F_main_BB_for_body_i_3 = 5'd3;
parameter [4:0] LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4 = 5'd4;
parameter [4:0] LEGUP_F_main_BB_for_cond10_preheader_i_5 = 5'd5;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_6 = 5'd6;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_7 = 5'd7;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_8 = 5'd8;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_9 = 5'd9;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_10 = 5'd10;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_11 = 5'd11;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_12 = 5'd12;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_13 = 5'd13;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_14 = 5'd14;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_15 = 5'd15;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_16 = 5'd16;
parameter [4:0] LEGUP_F_main_BB_for_body13_i_17 = 5'd17;
parameter [4:0] LEGUP_F_main_BB_for_inc74_i_18 = 5'd18;
parameter [4:0] LEGUP_F_main_BB_poly5_exit_19 = 5'd19;
parameter [4:0] LEGUP_F_main_BB_poly5_exit_20 = 5'd20;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [4:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [4:0] next_state;
wire  fsm_stall;
reg [10:0] main_for_body_i_k_0110_i;
reg [10:0] main_for_body_i_k_0110_i_reg;
reg [15:0] main_for_body_i_bit_select12;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx2_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx4_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx5_i;
reg [11:0] main_for_body_i_0;
reg [11:0] main_for_body_i_0_reg;
reg  main_for_body_i_exitcond5;
reg  main_for_body_i_exitcond5_reg;
reg [6:0] main_for_cond10_preheader_i_i_0109_i;
reg [6:0] main_for_cond10_preheader_i_i_0109_i_reg;
reg [31:0] main_for_body13_i_k_1108_i;
reg [31:0] main_for_body13_i_k_1108_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx14_i;
reg [31:0] main_for_body13_i_1;
reg [31:0] main_for_body13_i_1_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx18_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx22_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx41_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx70_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body13_i_arrayidx70_i_reg;
reg [15:0] main_for_body13_i_2;
reg [15:0] main_for_body13_i_2_reg;
reg [11:0] main_for_body13_i_bit_select8;
reg [9:0] main_for_body13_i_bit_select6;
reg [10:0] main_for_body13_i_bit_select4;
reg [7:0] main_for_body13_i_bit_select2;
reg [14:0] main_for_body13_i_bit_select;
reg [15:0] main_for_body13_i_3;
reg [15:0] main_for_body13_i_mul_i;
reg [15:0] main_for_body13_i_add_i;
reg [15:0] main_for_body13_i_mul20_i;
reg [15:0] main_for_body13_i_sub21_i;
reg [15:0] main_for_body13_i_4;
reg [15:0] main_for_body13_i_sr_negate;
reg [14:0] main_for_body13_i_bit_select10;
reg [15:0] main_for_body13_i_bit_concat11;
reg [15:0] main_for_body13_i_bit_concat9;
reg [15:0] main_for_body13_i_bit_concat7;
reg [15:0] main_for_body13_i_sr_add;
reg [15:0] main_for_body13_i_newEarly_sub30_i;
reg [15:0] main_for_body13_i_newCurOp_sub30_i;
reg [15:0] main_for_body13_i_mul31_i;
reg [15:0] main_for_body13_i_bit_concat5;
reg [15:0] main_for_body13_i_bit_concat3;
reg [15:0] main_for_body13_i_sr_add9;
reg [15:0] main_for_body13_i_sub37_i;
reg [15:0] main_for_body13_i_mul38_i;
reg [15:0] main_for_body13_i_add39_i;
reg [15:0] main_for_body13_i_add39_i_reg;
reg [15:0] main_for_body13_i_mul40_i;
reg [15:0] main_for_body13_i_5;
reg [15:0] main_for_body13_i_5_reg;
reg [15:0] main_for_body13_i_sub50_i;
reg [15:0] main_for_body13_i_mul51_i;
reg [15:0] main_for_body13_i_add52_i;
reg [15:0] main_for_body13_i_bit_concat1;
reg [15:0] main_for_body13_i_sub60_i;
reg [15:0] main_for_body13_i_add61_i;
reg [15:0] main_for_body13_i_mul62_i;
reg [15:0] main_for_body13_i_sub63_i;
reg [15:0] main_for_body13_i_mul64_i;
reg [15:0] main_for_body13_i_mul64_i_reg;
reg [15:0] main_for_body13_i_tmp_i;
reg [15:0] main_for_body13_i_tmp107_i;
reg [15:0] main_for_body13_i_tmp107_i_reg;
reg [15:0] main_for_body13_i_mul68_i;
reg [31:0] main_for_body13_i_6;
reg [31:0] main_for_body13_i_6_reg;
reg  main_for_body13_i_exitcond3;
reg  main_for_body13_i_exitcond3_reg;
reg [7:0] main_for_inc74_i_7;
reg  main_for_inc74_i_exitcond4;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_poly5_exit_arrayidx77_i;
reg [15:0] main_poly5_exit_8;
reg [31:0] main_poly5_exit_bit_concat;
reg [9:0] main_entry_a_i_address_a;
reg  main_entry_a_i_write_enable_a;
reg [15:0] main_entry_a_i_in_a;
wire [15:0] main_entry_a_i_out_a;
reg [9:0] main_entry_b_i_address_a;
reg  main_entry_b_i_write_enable_a;
reg [15:0] main_entry_b_i_in_a;
wire [15:0] main_entry_b_i_out_a;
reg [9:0] main_entry_c_i_address_a;
reg  main_entry_c_i_write_enable_a;
reg [15:0] main_entry_c_i_in_a;
wire [15:0] main_entry_c_i_out_a;
reg [9:0] main_entry_out_i_address_a;
reg  main_entry_out_i_write_enable_a;
reg [15:0] main_entry_out_i_in_a;
wire [15:0] main_entry_out_i_out_a;
reg [15:0] main_for_body_i_k_0110_i_reg_width_extended;
wire  main_for_body13_i_bit_concat11_bit_select_operand_2;
wire [3:0] main_for_body13_i_bit_concat9_bit_select_operand_2;
wire [5:0] main_for_body13_i_bit_concat7_bit_select_operand_2;
reg [15:0] op0_main_for_body13_i_newCurOp_sub30_i_reg;
reg [15:0] op1_main_for_body13_i_2_reg;
reg  legup_mult_main_for_body13_i_mul31_i_en;
reg [15:0] main_for_body13_i_mul31_i_stage0_reg;
wire [4:0] main_for_body13_i_bit_concat5_bit_select_operand_2;
wire [7:0] main_for_body13_i_bit_concat3_bit_select_operand_2;
reg [15:0] op0_main_for_body13_i_4_reg;
reg [15:0] op1_main_for_body13_i_sub37_i_reg;
reg  legup_mult_main_for_body13_i_mul38_i_en;
reg [15:0] main_for_body13_i_mul38_i_stage0_reg;
reg [15:0] op0_main_for_body13_i_sub50_i_reg;
reg  legup_mult_main_for_body13_i_mul51_i_en;
reg [15:0] main_for_body13_i_mul51_i_stage0_reg;
wire  main_for_body13_i_bit_concat1_bit_select_operand_2;
reg [15:0] op0_main_for_body13_i_add61_i_reg;
reg [15:0] op1_main_for_body13_i_4_reg;
reg  legup_mult_main_for_body13_i_mul62_i_en;
reg [15:0] main_for_body13_i_mul62_i_stage0_reg;
reg [15:0] op0_main_for_body13_i_5_reg;
reg  legup_mult_main_for_body13_i_tmp107_i_en;
reg [15:0] main_for_body13_i_tmp107_i_stage0_reg;
reg [15:0] op0_main_for_body13_i_3_reg;
reg [15:0] op1_main_for_body13_i_2_reg_reg;
reg  legup_mult_main_for_body13_i_mul_i_en;
reg [15:0] main_for_body13_i_mul_i_stage0_reg;
reg [15:0] op0_main_for_body13_i_sub63_i_reg;
reg [15:0] op1_main_for_body13_i_5_reg_reg;
reg  legup_mult_main_for_body13_i_mul64_i_en;
reg [15:0] main_for_body13_i_mul64_i_stage0_reg;
reg [15:0] op0_main_for_body13_i_add_i_reg;
reg  legup_mult_main_for_body13_i_mul20_i_en;
reg [15:0] main_for_body13_i_mul20_i_stage0_reg;
reg [15:0] op0_main_for_body13_i_sub21_i_reg;
reg [15:0] op1_main_for_body13_i_add39_i_reg_reg;
reg  legup_mult_main_for_body13_i_mul40_i_en;
reg [15:0] main_for_body13_i_mul40_i_stage0_reg;
reg [15:0] op0_main_for_body13_i_tmp107_i_reg_reg;
reg [15:0] op1_main_for_body13_i_tmp_i_reg;
reg  legup_mult_main_for_body13_i_mul68_i_en;
reg [15:0] main_for_body13_i_mul68_i_stage0_reg;
wire [15:0] main_poly5_exit_bit_concat_bit_select_operand_0;



//   %a.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port main_entry_a_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_a_i_address_a ),
	.wren_a( main_entry_a_i_write_enable_a ),
	.data_a( main_entry_a_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_a_i_out_a )
);
defparam main_entry_a_i.width_a = 16;
defparam main_entry_a_i.widthad_a = 10;
defparam main_entry_a_i.width_be_a = 2;
defparam main_entry_a_i.numwords_a = 1024;
defparam main_entry_a_i.latency = 1;


//   %b.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port main_entry_b_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_b_i_address_a ),
	.wren_a( main_entry_b_i_write_enable_a ),
	.data_a( main_entry_b_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_b_i_out_a )
);
defparam main_entry_b_i.width_a = 16;
defparam main_entry_b_i.widthad_a = 10;
defparam main_entry_b_i.width_be_a = 2;
defparam main_entry_b_i.numwords_a = 1024;
defparam main_entry_b_i.latency = 1;


//   %c.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port main_entry_c_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_c_i_address_a ),
	.wren_a( main_entry_c_i_write_enable_a ),
	.data_a( main_entry_c_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_c_i_out_a )
);
defparam main_entry_c_i.width_a = 16;
defparam main_entry_c_i.widthad_a = 10;
defparam main_entry_c_i.width_be_a = 2;
defparam main_entry_c_i.numwords_a = 1024;
defparam main_entry_c_i.latency = 1;


//   %out.i = alloca [1024 x i16], align 2, !dbg !31, !MSB !32, !LSB !33, !extendFrom !32
ram_single_port main_entry_out_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_out_i_address_a ),
	.wren_a( main_entry_out_i_write_enable_a ),
	.data_a( main_entry_out_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_out_i_out_a )
);
defparam main_entry_out_i.width_a = 16;
defparam main_entry_out_i.widthad_a = 10;
defparam main_entry_out_i.width_be_a = 2;
defparam main_entry_out_i.numwords_a = 1024;
defparam main_entry_out_i.latency = 1;

/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_poly5_exit_20)) begin
		$write("%d\n", $signed(main_poly5_exit_bit_concat));
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_for_body_i_2;
LEGUP_F_main_BB_for_body13_i_10:
		next_state = LEGUP_F_main_BB_for_body13_i_11;
LEGUP_F_main_BB_for_body13_i_11:
		next_state = LEGUP_F_main_BB_for_body13_i_12;
LEGUP_F_main_BB_for_body13_i_12:
		next_state = LEGUP_F_main_BB_for_body13_i_13;
LEGUP_F_main_BB_for_body13_i_13:
		next_state = LEGUP_F_main_BB_for_body13_i_14;
LEGUP_F_main_BB_for_body13_i_14:
		next_state = LEGUP_F_main_BB_for_body13_i_15;
LEGUP_F_main_BB_for_body13_i_15:
		next_state = LEGUP_F_main_BB_for_body13_i_16;
LEGUP_F_main_BB_for_body13_i_16:
		next_state = LEGUP_F_main_BB_for_body13_i_17;
LEGUP_F_main_BB_for_body13_i_17:
	if ((fsm_stall == 1'd0) && (main_for_body13_i_exitcond3_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc74_i_18;
	else if ((fsm_stall == 1'd0) && (main_for_body13_i_exitcond3_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body13_i_6;
LEGUP_F_main_BB_for_body13_i_6:
		next_state = LEGUP_F_main_BB_for_body13_i_7;
LEGUP_F_main_BB_for_body13_i_7:
		next_state = LEGUP_F_main_BB_for_body13_i_8;
LEGUP_F_main_BB_for_body13_i_8:
		next_state = LEGUP_F_main_BB_for_body13_i_9;
LEGUP_F_main_BB_for_body13_i_9:
		next_state = LEGUP_F_main_BB_for_body13_i_10;
LEGUP_F_main_BB_for_body_i_2:
		next_state = LEGUP_F_main_BB_for_body_i_3;
LEGUP_F_main_BB_for_body_i_3:
	if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond5_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond5_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_2;
LEGUP_F_main_BB_for_cond10_preheader_i_5:
		next_state = LEGUP_F_main_BB_for_body13_i_6;
LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4:
		next_state = LEGUP_F_main_BB_for_cond10_preheader_i_5;
LEGUP_F_main_BB_for_inc74_i_18:
	if ((fsm_stall == 1'd0) && (main_for_inc74_i_exitcond4 == 1'd1))
		next_state = LEGUP_F_main_BB_poly5_exit_19;
	else if ((fsm_stall == 1'd0) && (main_for_inc74_i_exitcond4 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond10_preheader_i_5;
LEGUP_F_main_BB_poly5_exit_19:
		next_state = LEGUP_F_main_BB_poly5_exit_20;
LEGUP_F_main_BB_poly5_exit_20:
		next_state = LEGUP_0;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_i_k_0110_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_i_3) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond5_reg == 1'd0))) */ begin
		main_for_body_i_k_0110_i = main_for_body_i_0_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_i_k_0110_i_reg <= main_for_body_i_k_0110_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_3) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond5_reg == 1'd0))) begin
		main_for_body_i_k_0110_i_reg <= main_for_body_i_k_0110_i;
	end
end
always @(*) begin
		main_for_body_i_bit_select12 = main_for_body_i_k_0110_i_reg_width_extended[15:0];
end
always @(*) begin
		main_for_body_i_arrayidx_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0110_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx2_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0110_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx4_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0110_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx5_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_0110_i_reg}));
end
always @(*) begin
		main_for_body_i_0 = ({1'd0,main_for_body_i_k_0110_i_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_for_body_i_0_reg <= main_for_body_i_0;
	end
end
always @(*) begin
		main_for_body_i_exitcond5 = (main_for_body_i_0 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_for_body_i_exitcond5_reg <= main_for_body_i_exitcond5;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_cond10_preheader_i_i_0109_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc74_i_18) & (fsm_stall == 1'd0)) & (main_for_inc74_i_exitcond4 == 1'd0))) */ begin
		main_for_cond10_preheader_i_i_0109_i = main_for_inc74_i_7;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_cond10_preheader_i_i_0109_i_reg <= main_for_cond10_preheader_i_i_0109_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc74_i_18) & (fsm_stall == 1'd0)) & (main_for_inc74_i_exitcond4 == 1'd0))) begin
		main_for_cond10_preheader_i_i_0109_i_reg <= main_for_cond10_preheader_i_i_0109_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_5) & (fsm_stall == 1'd0))) begin
		main_for_body13_i_k_1108_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body13_i_17) & (fsm_stall == 1'd0)) & (main_for_body13_i_exitcond3_reg == 1'd0))) */ begin
		main_for_body13_i_k_1108_i = main_for_body13_i_6_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond10_preheader_i_5) & (fsm_stall == 1'd0))) begin
		main_for_body13_i_k_1108_i_reg <= main_for_body13_i_k_1108_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body13_i_17) & (fsm_stall == 1'd0)) & (main_for_body13_i_exitcond3_reg == 1'd0))) begin
		main_for_body13_i_k_1108_i_reg <= main_for_body13_i_k_1108_i;
	end
end
always @(*) begin
		main_for_body13_i_arrayidx14_i = (1'd0 + (2 * main_for_body13_i_k_1108_i_reg));
end
always @(*) begin
		main_for_body13_i_1 = (main_for_body13_i_k_1108_i_reg + $signed(-32'd432));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_for_body13_i_1_reg <= main_for_body13_i_1;
	end
end
always @(*) begin
		main_for_body13_i_arrayidx18_i = (1'd0 + (2 * main_for_body13_i_1_reg));
end
always @(*) begin
		main_for_body13_i_arrayidx22_i = (1'd0 + (2 * main_for_body13_i_k_1108_i_reg));
end
always @(*) begin
		main_for_body13_i_arrayidx41_i = (1'd0 + (2 * main_for_body13_i_k_1108_i_reg));
end
always @(*) begin
		main_for_body13_i_arrayidx70_i = (1'd0 + (2 * main_for_body13_i_k_1108_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_for_body13_i_arrayidx70_i_reg <= main_for_body13_i_arrayidx70_i;
	end
end
always @(*) begin
		main_for_body13_i_2 = main_entry_a_i_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_2_reg <= main_for_body13_i_2;
	end
end
always @(*) begin
		main_for_body13_i_bit_select8 = main_for_body13_i_2[11:0];
end
always @(*) begin
		main_for_body13_i_bit_select6 = main_for_body13_i_2[9:0];
end
always @(*) begin
		main_for_body13_i_bit_select4 = main_for_body13_i_2[10:0];
end
always @(*) begin
		main_for_body13_i_bit_select2 = main_for_body13_i_2[7:0];
end
always @(*) begin
		main_for_body13_i_bit_select = main_for_body13_i_2[14:0];
end
always @(*) begin
		main_for_body13_i_3 = main_entry_a_i_out_a;
end
always @(*) begin
	main_for_body13_i_mul_i = main_for_body13_i_mul_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_add_i = (main_for_body13_i_mul_i + $signed(-16'd3328));
end
always @(*) begin
	main_for_body13_i_mul20_i = main_for_body13_i_mul20_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sub21_i = (main_for_body13_i_mul20_i + 16'd28672);
end
always @(*) begin
		main_for_body13_i_4 = main_entry_b_i_out_a;
end
always @(*) begin
		main_for_body13_i_sr_negate = (16'd0 - main_for_body13_i_2);
end
always @(*) begin
		main_for_body13_i_bit_select10 = main_for_body13_i_sr_negate[14:0];
end
always @(*) begin
		main_for_body13_i_bit_concat11 = {main_for_body13_i_bit_select10[14:0], main_for_body13_i_bit_concat11_bit_select_operand_2};
end
always @(*) begin
		main_for_body13_i_bit_concat9 = {main_for_body13_i_bit_select8[11:0], main_for_body13_i_bit_concat9_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body13_i_bit_concat7 = {main_for_body13_i_bit_select6[9:0], main_for_body13_i_bit_concat7_bit_select_operand_2[5:0]};
end
always @(*) begin
		main_for_body13_i_sr_add = (main_for_body13_i_bit_concat11 + main_for_body13_i_bit_concat9);
end
always @(*) begin
		main_for_body13_i_newEarly_sub30_i = (main_for_body13_i_bit_concat7 + -16'd9504);
end
always @(*) begin
		main_for_body13_i_newCurOp_sub30_i = (main_for_body13_i_newEarly_sub30_i + main_for_body13_i_sr_add);
end
always @(*) begin
	main_for_body13_i_mul31_i = main_for_body13_i_mul31_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_bit_concat5 = {main_for_body13_i_bit_select4[10:0], main_for_body13_i_bit_concat5_bit_select_operand_2[4:0]};
end
always @(*) begin
		main_for_body13_i_bit_concat3 = {main_for_body13_i_bit_select2[7:0], main_for_body13_i_bit_concat3_bit_select_operand_2[7:0]};
end
always @(*) begin
		main_for_body13_i_sr_add9 = (main_for_body13_i_bit_concat5 + main_for_body13_i_bit_concat3);
end
always @(*) begin
		main_for_body13_i_sub37_i = (main_for_body13_i_sr_add9 + $signed(-16'd5184));
end
always @(*) begin
	main_for_body13_i_mul38_i = main_for_body13_i_mul38_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_add39_i = (main_for_body13_i_mul31_i + main_for_body13_i_mul38_i);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_9)) begin
		main_for_body13_i_add39_i_reg <= main_for_body13_i_add39_i;
	end
end
always @(*) begin
	main_for_body13_i_mul40_i = main_for_body13_i_mul40_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_5 = main_entry_c_i_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_for_body13_i_5_reg <= main_for_body13_i_5;
	end
end
always @(*) begin
		main_for_body13_i_sub50_i = (main_for_body13_i_2 + $signed(-16'd207));
end
always @(*) begin
	main_for_body13_i_mul51_i = main_for_body13_i_mul51_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_add52_i = (main_for_body13_i_mul51_i + 16'd3456);
end
always @(*) begin
		main_for_body13_i_bit_concat1 = {main_for_body13_i_bit_select[14:0], main_for_body13_i_bit_concat1_bit_select_operand_2};
end
always @(*) begin
		main_for_body13_i_sub60_i = (main_for_body13_i_bit_concat1 + 16'd144);
end
always @(*) begin
		main_for_body13_i_add61_i = (main_for_body13_i_sub60_i - main_for_body13_i_5);
end
always @(*) begin
	main_for_body13_i_mul62_i = main_for_body13_i_mul62_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_sub63_i = (main_for_body13_i_add52_i - main_for_body13_i_mul62_i);
end
always @(*) begin
	main_for_body13_i_mul64_i = main_for_body13_i_mul64_i_stage0_reg;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_11)) begin
		main_for_body13_i_mul64_i_reg <= main_for_body13_i_mul64_i;
	end
end
always @(*) begin
		main_for_body13_i_tmp_i = (main_for_body13_i_mul64_i_reg + main_for_body13_i_mul40_i);
end
always @(*) begin
	main_for_body13_i_tmp107_i = main_for_body13_i_tmp107_i_stage0_reg;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_9)) begin
		main_for_body13_i_tmp107_i_reg <= main_for_body13_i_tmp107_i;
	end
end
always @(*) begin
	main_for_body13_i_mul68_i = main_for_body13_i_mul68_i_stage0_reg;
end
always @(*) begin
		main_for_body13_i_6 = (main_for_body13_i_k_1108_i_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_for_body13_i_6_reg <= main_for_body13_i_6;
	end
end
always @(*) begin
		main_for_body13_i_exitcond3 = (main_for_body13_i_6 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_for_body13_i_exitcond3_reg <= main_for_body13_i_exitcond3;
	end
end
always @(*) begin
		main_for_inc74_i_7 = ({1'd0,main_for_cond10_preheader_i_i_0109_i_reg} + 32'd1);
end
always @(*) begin
		main_for_inc74_i_exitcond4 = (main_for_inc74_i_7 == 32'd100);
end
assign main_poly5_exit_arrayidx77_i = (1'd0 + (2 * 32'd50));
always @(*) begin
		main_poly5_exit_8 = main_entry_out_i_out_a;
end
always @(*) begin
		main_poly5_exit_bit_concat = {main_poly5_exit_bit_concat_bit_select_operand_0[15:0], main_poly5_exit_8[15:0]};
end
always @(*) begin
	main_entry_a_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_a_i_address_a = (main_for_body_i_arrayidx_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_entry_a_i_address_a = (main_for_body13_i_arrayidx14_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		main_entry_a_i_address_a = (main_for_body13_i_arrayidx18_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_a_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_a_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_a_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_a_i_in_a = main_for_body_i_bit_select12;
	end
end
always @(*) begin
	main_entry_b_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_b_i_address_a = (main_for_body_i_arrayidx2_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_entry_b_i_address_a = (main_for_body13_i_arrayidx22_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_b_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_b_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_b_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_b_i_in_a = main_for_body_i_bit_select12;
	end
end
always @(*) begin
	main_entry_c_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_c_i_address_a = (main_for_body_i_arrayidx4_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_6)) begin
		main_entry_c_i_address_a = (main_for_body13_i_arrayidx41_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_c_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_c_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_c_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_c_i_in_a = main_for_body_i_bit_select12;
	end
end
always @(*) begin
	main_entry_out_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_out_i_address_a = (main_for_body_i_arrayidx5_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_16)) begin
		main_entry_out_i_address_a = (main_for_body13_i_arrayidx70_i_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_poly5_exit_19)) begin
		main_entry_out_i_address_a = (main_poly5_exit_arrayidx77_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_out_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_out_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_16)) begin
		main_entry_out_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_out_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_out_i_in_a = 16'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_16)) begin
		main_entry_out_i_in_a = main_for_body13_i_mul68_i;
	end
end
always @(*) begin
	main_for_body_i_k_0110_i_reg_width_extended = {5'd0,main_for_body_i_k_0110_i_reg};
end
assign main_for_body13_i_bit_concat11_bit_select_operand_2 = 1'd0;
assign main_for_body13_i_bit_concat9_bit_select_operand_2 = 4'd0;
assign main_for_body13_i_bit_concat7_bit_select_operand_2 = 6'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op0_main_for_body13_i_newCurOp_sub30_i_reg <= main_for_body13_i_newCurOp_sub30_i;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op1_main_for_body13_i_2_reg <= main_for_body13_i_2;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op1_main_for_body13_i_2_reg <= main_for_body13_i_2;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul31_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul31_i_en == 1'd1)) begin
		main_for_body13_i_mul31_i_stage0_reg <= (op0_main_for_body13_i_newCurOp_sub30_i_reg * op1_main_for_body13_i_2_reg);
	end
end
assign main_for_body13_i_bit_concat5_bit_select_operand_2 = 5'd0;
assign main_for_body13_i_bit_concat3_bit_select_operand_2 = 8'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op0_main_for_body13_i_4_reg <= main_for_body13_i_4;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op1_main_for_body13_i_sub37_i_reg <= main_for_body13_i_sub37_i;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul38_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul38_i_en == 1'd1)) begin
		main_for_body13_i_mul38_i_stage0_reg <= (op0_main_for_body13_i_4_reg * op1_main_for_body13_i_sub37_i_reg);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op0_main_for_body13_i_sub50_i_reg <= main_for_body13_i_sub50_i;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul51_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul51_i_en == 1'd1)) begin
		main_for_body13_i_mul51_i_stage0_reg <= (op0_main_for_body13_i_sub50_i_reg * op1_main_for_body13_i_2_reg);
	end
end
assign main_for_body13_i_bit_concat1_bit_select_operand_2 = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op0_main_for_body13_i_add61_i_reg <= main_for_body13_i_add61_i;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op1_main_for_body13_i_4_reg <= main_for_body13_i_4;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op1_main_for_body13_i_4_reg <= main_for_body13_i_4;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul62_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul62_i_en == 1'd1)) begin
		main_for_body13_i_mul62_i_stage0_reg <= (op0_main_for_body13_i_add61_i_reg * op1_main_for_body13_i_4_reg);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_7)) begin
		op0_main_for_body13_i_5_reg <= main_for_body13_i_5;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_tmp107_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_tmp107_i_en == 1'd1)) begin
		main_for_body13_i_tmp107_i_stage0_reg <= (op0_main_for_body13_i_5_reg * op1_main_for_body13_i_4_reg);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_8)) begin
		op0_main_for_body13_i_3_reg <= main_for_body13_i_3;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_8)) begin
		op1_main_for_body13_i_2_reg_reg <= main_for_body13_i_2_reg;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_10)) begin
		op1_main_for_body13_i_2_reg_reg <= main_for_body13_i_2_reg;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul_i_en == 1'd1)) begin
		main_for_body13_i_mul_i_stage0_reg <= (op0_main_for_body13_i_3_reg * op1_main_for_body13_i_2_reg_reg);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_9)) begin
		op0_main_for_body13_i_sub63_i_reg <= main_for_body13_i_sub63_i;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_9)) begin
		op1_main_for_body13_i_5_reg_reg <= main_for_body13_i_5_reg;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul64_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul64_i_en == 1'd1)) begin
		main_for_body13_i_mul64_i_stage0_reg <= (op0_main_for_body13_i_sub63_i_reg * op1_main_for_body13_i_5_reg_reg);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_10)) begin
		op0_main_for_body13_i_add_i_reg <= main_for_body13_i_add_i;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul20_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul20_i_en == 1'd1)) begin
		main_for_body13_i_mul20_i_stage0_reg <= (op0_main_for_body13_i_add_i_reg * op1_main_for_body13_i_2_reg_reg);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_12)) begin
		op0_main_for_body13_i_sub21_i_reg <= main_for_body13_i_sub21_i;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_12)) begin
		op1_main_for_body13_i_add39_i_reg_reg <= main_for_body13_i_add39_i_reg;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul40_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul40_i_en == 1'd1)) begin
		main_for_body13_i_mul40_i_stage0_reg <= (op0_main_for_body13_i_sub21_i_reg * op1_main_for_body13_i_add39_i_reg_reg);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_14)) begin
		op0_main_for_body13_i_tmp107_i_reg_reg <= main_for_body13_i_tmp107_i_reg;
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body13_i_14)) begin
		op1_main_for_body13_i_tmp_i_reg <= main_for_body13_i_tmp_i;
	end
end
always @(*) begin
	legup_mult_main_for_body13_i_mul68_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body13_i_mul68_i_en == 1'd1)) begin
		main_for_body13_i_mul68_i_stage0_reg <= (op0_main_for_body13_i_tmp107_i_reg_reg * op1_main_for_body13_i_tmp_i_reg);
	end
end
assign main_poly5_exit_bit_concat_bit_select_operand_0 = 16'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_poly5_exit_20)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_poly5_exit_20)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a,
	address_b,
	wren_b,
	data_b,
	byteena_b,
	q_b
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_be_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  width_be_b = 1'd0;
parameter  init_file_mem = {`MEM_INIT_DIR, "UNUSED.mem"};
parameter  latency = 1;

input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
reg [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
reg [(width_b-1):0] q_b_wire;
input  wren_b;
input [(width_a-1):0] data_b;
input [width_be_a-1:0] byteena_b;

reg [width_a-1:0] ram [numwords_a-1:0];

initial begin
	if (init_file_mem != {`MEM_INIT_DIR, "UNUSED.mem"})
        $readmemb(init_file_mem, ram);
end

localparam input_latency = ((latency - 1) >> 1);
localparam output_latency = (latency - 1) - input_latency;
integer j;

reg [(widthad_a-1):0] address_a_reg[input_latency:0];
reg  wren_a_reg[input_latency:0];
reg [(width_a-1):0] data_a_reg[input_latency:0];
reg [(width_be_a-1):0] byteena_a_reg[input_latency:0];
reg [(widthad_b-1):0] address_b_reg[input_latency:0];
reg  wren_b_reg[input_latency:0];
reg [(width_b-1):0] data_b_reg[input_latency:0];
reg [(width_be_b-1):0] byteena_b_reg[input_latency:0];

always @(*)
begin
  address_a_reg[0] = address_a;
  wren_a_reg[0] = wren_a;
  data_a_reg[0] = data_a;
  byteena_a_reg[0] = byteena_a;
  address_b_reg[0] = address_b;
  wren_b_reg[0] = wren_b;
  data_b_reg[0] = data_b;
  byteena_b_reg[0] = byteena_b;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < input_latency; j=j+1)
   begin
       address_a_reg[j+1] <= address_a_reg[j];
       wren_a_reg[j+1] <= wren_a_reg[j];
       data_a_reg[j+1] <= data_a_reg[j];
       byteena_a_reg[j+1] <= byteena_a_reg[j];
       address_b_reg[j+1] <= address_b_reg[j];
       wren_b_reg[j+1] <= wren_b_reg[j];
       data_b_reg[j+1] <= data_b_reg[j];
       byteena_b_reg[j+1] <= byteena_b_reg[j];
   end
end

always @ (posedge clk)
begin
    if (clken)
    begin // Port a
        if (wren_a_reg[input_latency])
        begin
            ram[address_a_reg[input_latency]] <= data_a_reg[input_latency];
            q_a_wire <= data_a_reg[input_latency];
        end
        else begin
            q_a_wire <= ram[address_a_reg[input_latency]];
        end
    end
end

always @ (posedge clk)
begin
    if (clken)
    begin // Port b
        if (wren_b_reg[input_latency])
        begin
            ram[address_b_reg[input_latency]] <= data_b_reg[input_latency];
            q_b_wire <= data_b_reg[input_latency];
        end
        else begin
            q_b_wire <= ram[address_b_reg[input_latency]];
        end
    end
end


reg [(width_a-1):0] q_a_reg[output_latency:0];

always @(*)
begin
   q_a_reg[0] <= q_a_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_a_reg[j+1] <= q_a_reg[j];
   end
end

assign q_a = q_a_reg[output_latency];
reg [(width_b-1):0] q_b_reg[output_latency:0];

always @(*)
begin
   q_b_reg[0] <= q_b_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_b_reg[j+1] <= q_b_reg[j];
   end
end

assign q_b = q_b_reg[output_latency];

endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
