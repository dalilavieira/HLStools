module emscripten_compute_dom_pk_code (
		input  wire        clock,                       //                       clock.clk
		input  wire        resetn,                      //                       reset.reset_n
		input  wire        start,                       //                        call.valid
		output wire        busy,                        //                            .stall
		output wire        done,                        //                      return.valid
		input  wire        stall,                       //                            .stall
		output wire [31:0] returndata,                  //                  returndata.data
		input  wire [63:0] keyCodeString,               //               keyCodeString.data
		input  wire [63:0] DOM_PK_0,                    //                    DOM_PK_0.data
		input  wire [63:0] DOM_PK_1,                    //                    DOM_PK_1.data
		input  wire [63:0] DOM_PK_2,                    //                    DOM_PK_2.data
		input  wire [63:0] DOM_PK_3,                    //                    DOM_PK_3.data
		input  wire [63:0] DOM_PK_4,                    //                    DOM_PK_4.data
		input  wire [63:0] DOM_PK_5,                    //                    DOM_PK_5.data
		input  wire [63:0] DOM_PK_6,                    //                    DOM_PK_6.data
		input  wire [63:0] DOM_PK_7,                    //                    DOM_PK_7.data
		input  wire [63:0] DOM_PK_8,                    //                    DOM_PK_8.data
		input  wire [63:0] DOM_PK_9,                    //                    DOM_PK_9.data
		input  wire [63:0] DOM_PK_A,                    //                    DOM_PK_A.data
		input  wire [63:0] DOM_PK_ALT_LEFT,             //             DOM_PK_ALT_LEFT.data
		input  wire [63:0] DOM_PK_ALT_RIGHT,            //            DOM_PK_ALT_RIGHT.data
		input  wire [63:0] DOM_PK_ARROW_DOWN,           //           DOM_PK_ARROW_DOWN.data
		input  wire [63:0] DOM_PK_ARROW_LEFT,           //           DOM_PK_ARROW_LEFT.data
		input  wire [63:0] DOM_PK_ARROW_RIGHT,          //          DOM_PK_ARROW_RIGHT.data
		input  wire [63:0] DOM_PK_ARROW_UP,             //             DOM_PK_ARROW_UP.data
		input  wire [63:0] DOM_PK_AUDIO_VOLUME_DOWN,    //    DOM_PK_AUDIO_VOLUME_DOWN.data
		input  wire [63:0] DOM_PK_AUDIO_VOLUME_MUTE,    //    DOM_PK_AUDIO_VOLUME_MUTE.data
		input  wire [63:0] DOM_PK_AUDIO_VOLUME_UP,      //      DOM_PK_AUDIO_VOLUME_UP.data
		input  wire [63:0] DOM_PK_B,                    //                    DOM_PK_B.data
		input  wire [63:0] DOM_PK_BACKQUOTE,            //            DOM_PK_BACKQUOTE.data
		input  wire [63:0] DOM_PK_BACKSLASH,            //            DOM_PK_BACKSLASH.data
		input  wire [63:0] DOM_PK_BACKSPACE,            //            DOM_PK_BACKSPACE.data
		input  wire [63:0] DOM_PK_BRACKET_LEFT,         //         DOM_PK_BRACKET_LEFT.data
		input  wire [63:0] DOM_PK_BRACKET_RIGHT,        //        DOM_PK_BRACKET_RIGHT.data
		input  wire [63:0] DOM_PK_BROWSER_BACK,         //         DOM_PK_BROWSER_BACK.data
		input  wire [63:0] DOM_PK_BROWSER_FAVORITES,    //    DOM_PK_BROWSER_FAVORITES.data
		input  wire [63:0] DOM_PK_BROWSER_FORWARD,      //      DOM_PK_BROWSER_FORWARD.data
		input  wire [63:0] DOM_PK_BROWSER_HOME,         //         DOM_PK_BROWSER_HOME.data
		input  wire [63:0] DOM_PK_BROWSER_REFRESH,      //      DOM_PK_BROWSER_REFRESH.data
		input  wire [63:0] DOM_PK_BROWSER_SEARCH,       //       DOM_PK_BROWSER_SEARCH.data
		input  wire [63:0] DOM_PK_BROWSER_STOP,         //         DOM_PK_BROWSER_STOP.data
		input  wire [63:0] DOM_PK_C,                    //                    DOM_PK_C.data
		input  wire [63:0] DOM_PK_CAPS_LOCK,            //            DOM_PK_CAPS_LOCK.data
		input  wire [63:0] DOM_PK_COMMA,                //                DOM_PK_COMMA.data
		input  wire [63:0] DOM_PK_CONTEXT_MENU,         //         DOM_PK_CONTEXT_MENU.data
		input  wire [63:0] DOM_PK_CONTROL_LEFT,         //         DOM_PK_CONTROL_LEFT.data
		input  wire [63:0] DOM_PK_CONTROL_RIGHT,        //        DOM_PK_CONTROL_RIGHT.data
		input  wire [63:0] DOM_PK_CONVERT,              //              DOM_PK_CONVERT.data
		input  wire [63:0] DOM_PK_COPY,                 //                 DOM_PK_COPY.data
		input  wire [63:0] DOM_PK_CUT,                  //                  DOM_PK_CUT.data
		input  wire [63:0] DOM_PK_D,                    //                    DOM_PK_D.data
		input  wire [63:0] DOM_PK_DELETE,               //               DOM_PK_DELETE.data
		input  wire [63:0] DOM_PK_E,                    //                    DOM_PK_E.data
		input  wire [63:0] DOM_PK_EJECT,                //                DOM_PK_EJECT.data
		input  wire [63:0] DOM_PK_END,                  //                  DOM_PK_END.data
		input  wire [63:0] DOM_PK_ENTER,                //                DOM_PK_ENTER.data
		input  wire [63:0] DOM_PK_EQUAL,                //                DOM_PK_EQUAL.data
		input  wire [63:0] DOM_PK_ESCAPE,               //               DOM_PK_ESCAPE.data
		input  wire [63:0] DOM_PK_F,                    //                    DOM_PK_F.data
		input  wire [63:0] DOM_PK_F1,                   //                   DOM_PK_F1.data
		input  wire [63:0] DOM_PK_F10,                  //                  DOM_PK_F10.data
		input  wire [63:0] DOM_PK_F11,                  //                  DOM_PK_F11.data
		input  wire [63:0] DOM_PK_F12,                  //                  DOM_PK_F12.data
		input  wire [63:0] DOM_PK_F13,                  //                  DOM_PK_F13.data
		input  wire [63:0] DOM_PK_F14,                  //                  DOM_PK_F14.data
		input  wire [63:0] DOM_PK_F15,                  //                  DOM_PK_F15.data
		input  wire [63:0] DOM_PK_F16,                  //                  DOM_PK_F16.data
		input  wire [63:0] DOM_PK_F17,                  //                  DOM_PK_F17.data
		input  wire [63:0] DOM_PK_F18,                  //                  DOM_PK_F18.data
		input  wire [63:0] DOM_PK_F19,                  //                  DOM_PK_F19.data
		input  wire [63:0] DOM_PK_F2,                   //                   DOM_PK_F2.data
		input  wire [63:0] DOM_PK_F20,                  //                  DOM_PK_F20.data
		input  wire [63:0] DOM_PK_F21,                  //                  DOM_PK_F21.data
		input  wire [63:0] DOM_PK_F22,                  //                  DOM_PK_F22.data
		input  wire [63:0] DOM_PK_F23,                  //                  DOM_PK_F23.data
		input  wire [63:0] DOM_PK_F24,                  //                  DOM_PK_F24.data
		input  wire [63:0] DOM_PK_F3,                   //                   DOM_PK_F3.data
		input  wire [63:0] DOM_PK_F4,                   //                   DOM_PK_F4.data
		input  wire [63:0] DOM_PK_F5,                   //                   DOM_PK_F5.data
		input  wire [63:0] DOM_PK_F6,                   //                   DOM_PK_F6.data
		input  wire [63:0] DOM_PK_F7,                   //                   DOM_PK_F7.data
		input  wire [63:0] DOM_PK_F8,                   //                   DOM_PK_F8.data
		input  wire [63:0] DOM_PK_F9,                   //                   DOM_PK_F9.data
		input  wire [63:0] DOM_PK_G,                    //                    DOM_PK_G.data
		input  wire [63:0] DOM_PK_H,                    //                    DOM_PK_H.data
		input  wire [63:0] DOM_PK_HELP,                 //                 DOM_PK_HELP.data
		input  wire [63:0] DOM_PK_HOME,                 //                 DOM_PK_HOME.data
		input  wire [63:0] DOM_PK_I,                    //                    DOM_PK_I.data
		input  wire [63:0] DOM_PK_INSERT,               //               DOM_PK_INSERT.data
		input  wire [63:0] DOM_PK_INTL_BACKSLASH,       //       DOM_PK_INTL_BACKSLASH.data
		input  wire [63:0] DOM_PK_INTL_RO,              //              DOM_PK_INTL_RO.data
		input  wire [63:0] DOM_PK_INTL_YEN,             //             DOM_PK_INTL_YEN.data
		input  wire [63:0] DOM_PK_J,                    //                    DOM_PK_J.data
		input  wire [63:0] DOM_PK_K,                    //                    DOM_PK_K.data
		input  wire [63:0] DOM_PK_KANA_MODE,            //            DOM_PK_KANA_MODE.data
		input  wire [63:0] DOM_PK_L,                    //                    DOM_PK_L.data
		input  wire [63:0] DOM_PK_LANG_1,               //               DOM_PK_LANG_1.data
		input  wire [63:0] DOM_PK_LANG_2,               //               DOM_PK_LANG_2.data
		input  wire [63:0] DOM_PK_LAUNCH_APP_1,         //         DOM_PK_LAUNCH_APP_1.data
		input  wire [63:0] DOM_PK_LAUNCH_APP_2,         //         DOM_PK_LAUNCH_APP_2.data
		input  wire [63:0] DOM_PK_LAUNCH_MAIL,          //          DOM_PK_LAUNCH_MAIL.data
		input  wire [63:0] DOM_PK_LAUNCH_MEDIA_PLAYER,  //  DOM_PK_LAUNCH_MEDIA_PLAYER.data
		input  wire [63:0] DOM_PK_M,                    //                    DOM_PK_M.data
		input  wire [63:0] DOM_PK_MEDIA_PLAY_PAUSE,     //     DOM_PK_MEDIA_PLAY_PAUSE.data
		input  wire [63:0] DOM_PK_MEDIA_SELECT,         //         DOM_PK_MEDIA_SELECT.data
		input  wire [63:0] DOM_PK_MEDIA_STOP,           //           DOM_PK_MEDIA_STOP.data
		input  wire [63:0] DOM_PK_MEDIA_TRACK_NEXT,     //     DOM_PK_MEDIA_TRACK_NEXT.data
		input  wire [63:0] DOM_PK_MEDIA_TRACK_PREVIOUS, // DOM_PK_MEDIA_TRACK_PREVIOUS.data
		input  wire [63:0] DOM_PK_META_LEFT,            //            DOM_PK_META_LEFT.data
		input  wire [63:0] DOM_PK_META_RIGHT,           //           DOM_PK_META_RIGHT.data
		input  wire [63:0] DOM_PK_MINUS,                //                DOM_PK_MINUS.data
		input  wire [63:0] DOM_PK_N,                    //                    DOM_PK_N.data
		input  wire [63:0] DOM_PK_NON_CONVERT,          //          DOM_PK_NON_CONVERT.data
		input  wire [63:0] DOM_PK_NUMPAD_0,             //             DOM_PK_NUMPAD_0.data
		input  wire [63:0] DOM_PK_NUMPAD_1,             //             DOM_PK_NUMPAD_1.data
		input  wire [63:0] DOM_PK_NUMPAD_2,             //             DOM_PK_NUMPAD_2.data
		input  wire [63:0] DOM_PK_NUMPAD_3,             //             DOM_PK_NUMPAD_3.data
		input  wire [63:0] DOM_PK_NUMPAD_4,             //             DOM_PK_NUMPAD_4.data
		input  wire [63:0] DOM_PK_NUMPAD_5,             //             DOM_PK_NUMPAD_5.data
		input  wire [63:0] DOM_PK_NUMPAD_6,             //             DOM_PK_NUMPAD_6.data
		input  wire [63:0] DOM_PK_NUMPAD_7,             //             DOM_PK_NUMPAD_7.data
		input  wire [63:0] DOM_PK_NUMPAD_8,             //             DOM_PK_NUMPAD_8.data
		input  wire [63:0] DOM_PK_NUMPAD_9,             //             DOM_PK_NUMPAD_9.data
		input  wire [63:0] DOM_PK_NUMPAD_ADD,           //           DOM_PK_NUMPAD_ADD.data
		input  wire [63:0] DOM_PK_NUMPAD_COMMA,         //         DOM_PK_NUMPAD_COMMA.data
		input  wire [63:0] DOM_PK_NUMPAD_DECIMAL,       //       DOM_PK_NUMPAD_DECIMAL.data
		input  wire [63:0] DOM_PK_NUMPAD_DIVIDE,        //        DOM_PK_NUMPAD_DIVIDE.data
		input  wire [63:0] DOM_PK_NUMPAD_ENTER,         //         DOM_PK_NUMPAD_ENTER.data
		input  wire [63:0] DOM_PK_NUMPAD_EQUAL,         //         DOM_PK_NUMPAD_EQUAL.data
		input  wire [63:0] DOM_PK_NUMPAD_MULTIPLY,      //      DOM_PK_NUMPAD_MULTIPLY.data
		input  wire [63:0] DOM_PK_NUMPAD_SUBTRACT,      //      DOM_PK_NUMPAD_SUBTRACT.data
		input  wire [63:0] DOM_PK_NUM_LOCK,             //             DOM_PK_NUM_LOCK.data
		input  wire [63:0] DOM_PK_O,                    //                    DOM_PK_O.data
		input  wire [63:0] DOM_PK_OS_LEFT,              //              DOM_PK_OS_LEFT.data
		input  wire [63:0] DOM_PK_OS_RIGHT,             //             DOM_PK_OS_RIGHT.data
		input  wire [63:0] DOM_PK_P,                    //                    DOM_PK_P.data
		input  wire [63:0] DOM_PK_PAGE_DOWN,            //            DOM_PK_PAGE_DOWN.data
		input  wire [63:0] DOM_PK_PAGE_UP,              //              DOM_PK_PAGE_UP.data
		input  wire [63:0] DOM_PK_PASTE,                //                DOM_PK_PASTE.data
		input  wire [63:0] DOM_PK_PAUSE,                //                DOM_PK_PAUSE.data
		input  wire [63:0] DOM_PK_PERIOD,               //               DOM_PK_PERIOD.data
		input  wire [63:0] DOM_PK_POWER,                //                DOM_PK_POWER.data
		input  wire [63:0] DOM_PK_PRINT_SCREEN,         //         DOM_PK_PRINT_SCREEN.data
		input  wire [63:0] DOM_PK_Q,                    //                    DOM_PK_Q.data
		input  wire [63:0] DOM_PK_QUOTE,                //                DOM_PK_QUOTE.data
		input  wire [63:0] DOM_PK_R,                    //                    DOM_PK_R.data
		input  wire [63:0] DOM_PK_S,                    //                    DOM_PK_S.data
		input  wire [63:0] DOM_PK_SCROLL_LOCK,          //          DOM_PK_SCROLL_LOCK.data
		input  wire [63:0] DOM_PK_SEMICOLON,            //            DOM_PK_SEMICOLON.data
		input  wire [63:0] DOM_PK_SHIFT_LEFT,           //           DOM_PK_SHIFT_LEFT.data
		input  wire [63:0] DOM_PK_SHIFT_RIGHT,          //          DOM_PK_SHIFT_RIGHT.data
		input  wire [63:0] DOM_PK_SLASH,                //                DOM_PK_SLASH.data
		input  wire [63:0] DOM_PK_SPACE,                //                DOM_PK_SPACE.data
		input  wire [63:0] DOM_PK_T,                    //                    DOM_PK_T.data
		input  wire [63:0] DOM_PK_TAB,                  //                  DOM_PK_TAB.data
		input  wire [63:0] DOM_PK_U,                    //                    DOM_PK_U.data
		input  wire [63:0] DOM_PK_UNKNOWN,              //              DOM_PK_UNKNOWN.data
		input  wire [63:0] DOM_PK_V,                    //                    DOM_PK_V.data
		input  wire [63:0] DOM_PK_W,                    //                    DOM_PK_W.data
		input  wire [63:0] DOM_PK_X,                    //                    DOM_PK_X.data
		input  wire [63:0] DOM_PK_Y,                    //                    DOM_PK_Y.data
		input  wire [63:0] DOM_PK_Z,                    //                    DOM_PK_Z.data
		output wire [63:0] avmm_0_rw_address,           //                   avmm_0_rw.address
		output wire [7:0]  avmm_0_rw_byteenable,        //                            .byteenable
		output wire        avmm_0_rw_read,              //                            .read
		input  wire [63:0] avmm_0_rw_readdata,          //                            .readdata
		output wire        avmm_0_rw_write,             //                            .write
		output wire [63:0] avmm_0_rw_writedata          //                            .writedata
	);
endmodule

