// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Mon Apr 20 09:42:08 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [4:0] LEGUP_0 = 5'd0;
parameter [4:0] LEGUP_F_main_BB_entry_1 = 5'd1;
parameter [4:0] LEGUP_F_main_BB_for_body_2 = 5'd2;
parameter [4:0] LEGUP_F_main_BB_for_body_3 = 5'd3;
parameter [4:0] LEGUP_F_main_BB_for_body_i_preheader_4 = 5'd4;
parameter [4:0] LEGUP_F_main_BB_for_inc32_us_i_5 = 5'd5;
parameter [4:0] LEGUP_F_main_BB_for_end27_us_us_i_6 = 5'd6;
parameter [4:0] LEGUP_F_main_BB_for_end27_us_us_i_7 = 5'd7;
parameter [4:0] LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8 = 5'd8;
parameter [4:0] LEGUP_F_main_BB_for_body15_us_us_i_9 = 5'd9;
parameter [4:0] LEGUP_F_main_BB_for_body15_us_us_i_10 = 5'd10;
parameter [4:0] LEGUP_F_main_BB_for_body15_us_us_i_11 = 5'd11;
parameter [4:0] LEGUP_F_main_BB_for_body15_us_us_i_12 = 5'd12;
parameter [4:0] LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_13 = 5'd13;
parameter [4:0] LEGUP_F_main_BB_for_body_i_14 = 5'd14;
parameter [4:0] LEGUP_F_main_BB_for_body_i_15 = 5'd15;
parameter [4:0] LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_preheader_16 = 5'd16;
parameter [4:0] LEGUP_F_main_BB_fir_exit_17 = 5'd17;
parameter [4:0] LEGUP_F_main_BB_fir_exit_18 = 5'd18;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [4:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [4:0] next_state;
wire  fsm_stall;
reg [5:0] main_for_body_k_05;
reg [5:0] main_for_body_k_05_reg;
reg [6:0] main_for_body_0;
reg [6:0] main_for_body_0_reg;
reg [15:0] main_for_body_bit_select1;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_arrayidx;
reg  main_for_body_exitcond4;
reg  main_for_body_exitcond4_reg;
reg [7:0] main_for_inc32_us_i_1;
reg  main_for_inc32_us_i_exitcond;
reg [31:0] main_for_end27_us_us_i_2;
reg [31:0] main_for_end27_us_us_i_2_reg;
reg  main_for_end27_us_us_i_exitcond2;
reg  main_for_end27_us_us_i_exitcond2_reg;
reg [31:0] main_for_body15_lr_ph_us_us_i_j_056_us_us_i;
reg [31:0] main_for_body15_lr_ph_us_us_i_j_056_us_us_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body15_lr_ph_us_us_i_arrayidx28_us_us_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body15_lr_ph_us_us_i_arrayidx28_us_us_i_reg;
reg [15:0] main_for_body15_us_us_i_fir_055_us_us_i;
reg [15:0] main_for_body15_us_us_i_fir_055_us_us_i_reg;
reg [31:0] main_for_body15_us_us_i_k_154_us_us_i;
reg [31:0] main_for_body15_us_us_i_k_154_us_us_i_reg;
reg [31:0] main_for_body15_us_us_i_3;
reg [31:0] main_for_body15_us_us_i_3_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body15_us_us_i_arrayidx17_us_us_i;
reg [31:0] main_for_body15_us_us_i_4;
reg [31:0] main_for_body15_us_us_i_4_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body15_us_us_i_arrayidx20_us_us_i;
reg [15:0] main_for_body15_us_us_i_5;
reg [15:0] main_for_body15_us_us_i_6;
reg [15:0] main_for_body15_us_us_i_mul_us_us_i;
reg [15:0] main_for_body15_us_us_i_add23_us_us_i;
reg [15:0] main_for_body15_us_us_i_add23_us_us_i_reg;
reg [31:0] main_for_body15_us_us_i_7;
reg [31:0] main_for_body15_us_us_i_7_reg;
reg  main_for_body15_us_us_i_exitcond1;
reg  main_for_body15_us_us_i_exitcond1_reg;
reg [6:0] main_for_cond8_preheader_split_us_us_i_i_058_us_i;
reg [6:0] main_for_cond8_preheader_split_us_us_i_i_058_us_i_reg;
reg [10:0] main_for_body_i_k_084_i;
reg [10:0] main_for_body_i_k_084_i_reg;
reg [15:0] main_for_body_i_bit_select;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx3_i;
reg [11:0] main_for_body_i_8;
reg [11:0] main_for_body_i_8_reg;
reg  main_for_body_i_exitcond3;
reg  main_for_body_i_exitcond3_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_fir_exit_arrayidx35_i;
reg [15:0] main_fir_exit_9;
reg [31:0] main_fir_exit_bit_concat;
reg [10:0] main_entry_vla_i1_address_a;
reg  main_entry_vla_i1_write_enable_a;
reg [15:0] main_entry_vla_i1_in_a;
wire [15:0] main_entry_vla_i1_out_a;
reg [10:0] main_entry_vla2_i2_address_a;
reg  main_entry_vla2_i2_write_enable_a;
reg [15:0] main_entry_vla2_i2_in_a;
wire [15:0] main_entry_vla2_i2_out_a;
reg [5:0] main_entry_coef_address_a;
reg  main_entry_coef_write_enable_a;
reg [15:0] main_entry_coef_in_a;
wire [15:0] main_entry_coef_out_a;
reg [15:0] main_for_body_0_width_extended;
reg  legup_mult_main_for_body15_us_us_i_mul_us_us_i_en;
reg [15:0] main_for_body15_us_us_i_mul_us_us_i_stage0_reg;
reg [15:0] main_for_body_i_k_084_i_reg_width_extended;
wire [15:0] main_fir_exit_bit_concat_bit_select_operand_0;



//   %vla.i1 = alloca [1087 x i16], align 2, !dbg !43, !MSB !45, !LSB !46, !extendFrom !45
ram_single_port_intel main_entry_vla_i1 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla_i1_address_a ),
	.wren_a( main_entry_vla_i1_write_enable_a ),
	.data_a( main_entry_vla_i1_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_vla_i1_out_a )
);
defparam main_entry_vla_i1.width_a = 16;
defparam main_entry_vla_i1.widthad_a = 11;
defparam main_entry_vla_i1.width_be_a = 2;
defparam main_entry_vla_i1.numwords_a = 1087;
defparam main_entry_vla_i1.latency = 1;


//   %vla2.i2 = alloca [1087 x i16], align 2, !dbg !47, !MSB !45, !LSB !46, !extendFrom !45
ram_single_port_intel main_entry_vla2_i2 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla2_i2_address_a ),
	.wren_a( main_entry_vla2_i2_write_enable_a ),
	.data_a( main_entry_vla2_i2_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_vla2_i2_out_a )
);
defparam main_entry_vla2_i2.width_a = 16;
defparam main_entry_vla2_i2.widthad_a = 11;
defparam main_entry_vla2_i2.width_be_a = 2;
defparam main_entry_vla2_i2.numwords_a = 1087;
defparam main_entry_vla2_i2.latency = 1;


//   %coef = alloca [63 x i16], align 2, !MSB !45, !LSB !46, !extendFrom !45
ram_single_port_intel main_entry_coef (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_coef_address_a ),
	.wren_a( main_entry_coef_write_enable_a ),
	.data_a( main_entry_coef_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_coef_out_a )
);
defparam main_entry_coef.width_a = 16;
defparam main_entry_coef.widthad_a = 6;
defparam main_entry_coef.width_be_a = 2;
defparam main_entry_coef.numwords_a = 63;
defparam main_entry_coef.latency = 1;

/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_fir_exit_18)) begin
		$write("%d\n", $signed(main_fir_exit_bit_concat));
		// to fix quartus warning
		if (reset == 1'b0 && ^(main_fir_exit_bit_concat) === 1'bX) finish <= 0;
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_for_body_2;
LEGUP_F_main_BB_fir_exit_17:
		next_state = LEGUP_F_main_BB_fir_exit_18;
LEGUP_F_main_BB_fir_exit_18:
		next_state = LEGUP_0;
LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8:
		next_state = LEGUP_F_main_BB_for_body15_us_us_i_9;
LEGUP_F_main_BB_for_body15_us_us_i_10:
		next_state = LEGUP_F_main_BB_for_body15_us_us_i_11;
LEGUP_F_main_BB_for_body15_us_us_i_11:
		next_state = LEGUP_F_main_BB_for_body15_us_us_i_12;
LEGUP_F_main_BB_for_body15_us_us_i_12:
	if ((fsm_stall == 1'd0) && (main_for_body15_us_us_i_exitcond1_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_end27_us_us_i_6;
	else if ((fsm_stall == 1'd0) && (main_for_body15_us_us_i_exitcond1_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body15_us_us_i_9;
LEGUP_F_main_BB_for_body15_us_us_i_9:
		next_state = LEGUP_F_main_BB_for_body15_us_us_i_10;
LEGUP_F_main_BB_for_body_2:
		next_state = LEGUP_F_main_BB_for_body_3;
LEGUP_F_main_BB_for_body_3:
	if ((fsm_stall == 1'd0) && (main_for_body_exitcond4_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_body_i_preheader_4;
	else if ((fsm_stall == 1'd0) && (main_for_body_exitcond4_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_2;
LEGUP_F_main_BB_for_body_i_14:
		next_state = LEGUP_F_main_BB_for_body_i_15;
LEGUP_F_main_BB_for_body_i_15:
	if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond3_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_preheader_16;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond3_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_14;
LEGUP_F_main_BB_for_body_i_preheader_4:
		next_state = LEGUP_F_main_BB_for_body_i_14;
LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_13:
		next_state = LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8;
LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_preheader_16:
		next_state = LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_13;
LEGUP_F_main_BB_for_end27_us_us_i_6:
		next_state = LEGUP_F_main_BB_for_end27_us_us_i_7;
LEGUP_F_main_BB_for_end27_us_us_i_7:
	if ((fsm_stall == 1'd0) && (main_for_end27_us_us_i_exitcond2_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc32_us_i_5;
	else if ((fsm_stall == 1'd0) && (main_for_end27_us_us_i_exitcond2_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8;
LEGUP_F_main_BB_for_inc32_us_i_5:
	if ((fsm_stall == 1'd0) && (main_for_inc32_us_i_exitcond == 1'd1))
		next_state = LEGUP_F_main_BB_fir_exit_17;
	else if ((fsm_stall == 1'd0) && (main_for_inc32_us_i_exitcond == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_13;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_k_05 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_3) & (fsm_stall == 1'd0)) & (main_for_body_exitcond4_reg == 1'd0))) */ begin
		main_for_body_k_05 = main_for_body_0_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_k_05_reg <= main_for_body_k_05;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_3) & (fsm_stall == 1'd0)) & (main_for_body_exitcond4_reg == 1'd0))) begin
		main_for_body_k_05_reg <= main_for_body_k_05;
	end
end
always @(*) begin
		main_for_body_0 = ({1'd0,main_for_body_k_05_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_for_body_0_reg <= main_for_body_0;
	end
end
always @(*) begin
		main_for_body_bit_select1 = main_for_body_0_width_extended[15:0];
end
always @(*) begin
		main_for_body_arrayidx = (1'd0 + (2 * {26'd0,main_for_body_k_05_reg}));
end
always @(*) begin
		main_for_body_exitcond4 = (main_for_body_0 == 32'd63);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_for_body_exitcond4_reg <= main_for_body_exitcond4;
	end
end
always @(*) begin
		main_for_inc32_us_i_1 = ({1'd0,main_for_cond8_preheader_split_us_us_i_i_058_us_i_reg} + 32'd1);
end
always @(*) begin
		main_for_inc32_us_i_exitcond = (main_for_inc32_us_i_1 == 32'd100);
end
always @(*) begin
		main_for_end27_us_us_i_2 = (main_for_body15_lr_ph_us_us_i_j_056_us_us_i_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_end27_us_us_i_6)) begin
		main_for_end27_us_us_i_2_reg <= main_for_end27_us_us_i_2;
	end
end
always @(*) begin
		main_for_end27_us_us_i_exitcond2 = (main_for_end27_us_us_i_2 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_end27_us_us_i_6)) begin
		main_for_end27_us_us_i_exitcond2_reg <= main_for_end27_us_us_i_exitcond2;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_end27_us_us_i_7) & (fsm_stall == 1'd0)) & (main_for_end27_us_us_i_exitcond2_reg == 1'd0))) begin
		main_for_body15_lr_ph_us_us_i_j_056_us_us_i = main_for_end27_us_us_i_2_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_13) & (fsm_stall == 1'd0))) */ begin
		main_for_body15_lr_ph_us_us_i_j_056_us_us_i = 32'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_end27_us_us_i_7) & (fsm_stall == 1'd0)) & (main_for_end27_us_us_i_exitcond2_reg == 1'd0))) begin
		main_for_body15_lr_ph_us_us_i_j_056_us_us_i_reg <= main_for_body15_lr_ph_us_us_i_j_056_us_us_i;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_13) & (fsm_stall == 1'd0))) begin
		main_for_body15_lr_ph_us_us_i_j_056_us_us_i_reg <= main_for_body15_lr_ph_us_us_i_j_056_us_us_i;
	end
end
always @(*) begin
		main_for_body15_lr_ph_us_us_i_arrayidx28_us_us_i = (1'd0 + (2 * main_for_body15_lr_ph_us_us_i_j_056_us_us_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8)) begin
		main_for_body15_lr_ph_us_us_i_arrayidx28_us_us_i_reg <= main_for_body15_lr_ph_us_us_i_arrayidx28_us_us_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8) & (fsm_stall == 1'd0))) begin
		main_for_body15_us_us_i_fir_055_us_us_i = 16'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_12) & (fsm_stall == 1'd0)) & (main_for_body15_us_us_i_exitcond1_reg == 1'd0))) */ begin
		main_for_body15_us_us_i_fir_055_us_us_i = main_for_body15_us_us_i_add23_us_us_i;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8) & (fsm_stall == 1'd0))) begin
		main_for_body15_us_us_i_fir_055_us_us_i_reg <= main_for_body15_us_us_i_fir_055_us_us_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_12) & (fsm_stall == 1'd0)) & (main_for_body15_us_us_i_exitcond1_reg == 1'd0))) begin
		main_for_body15_us_us_i_fir_055_us_us_i_reg <= main_for_body15_us_us_i_fir_055_us_us_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8) & (fsm_stall == 1'd0))) begin
		main_for_body15_us_us_i_k_154_us_us_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_12) & (fsm_stall == 1'd0)) & (main_for_body15_us_us_i_exitcond1_reg == 1'd0))) */ begin
		main_for_body15_us_us_i_k_154_us_us_i = main_for_body15_us_us_i_7_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body15_lr_ph_us_us_i_8) & (fsm_stall == 1'd0))) begin
		main_for_body15_us_us_i_k_154_us_us_i_reg <= main_for_body15_us_us_i_k_154_us_us_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_12) & (fsm_stall == 1'd0)) & (main_for_body15_us_us_i_exitcond1_reg == 1'd0))) begin
		main_for_body15_us_us_i_k_154_us_us_i_reg <= main_for_body15_us_us_i_k_154_us_us_i;
	end
end
always @(*) begin
		main_for_body15_us_us_i_3 = (main_for_body15_lr_ph_us_us_i_j_056_us_us_i_reg + main_for_body15_us_us_i_k_154_us_us_i_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_9)) begin
		main_for_body15_us_us_i_3_reg <= main_for_body15_us_us_i_3;
	end
end
always @(*) begin
		main_for_body15_us_us_i_arrayidx17_us_us_i = (1'd0 + (2 * main_for_body15_us_us_i_3_reg));
end
always @(*) begin
		main_for_body15_us_us_i_4 = (32'd62 - main_for_body15_us_us_i_k_154_us_us_i_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_9)) begin
		main_for_body15_us_us_i_4_reg <= main_for_body15_us_us_i_4;
	end
end
always @(*) begin
		main_for_body15_us_us_i_arrayidx20_us_us_i = (1'd0 + (2 * main_for_body15_us_us_i_4_reg));
end
always @(*) begin
		main_for_body15_us_us_i_5 = main_entry_vla_i1_out_a;
end
always @(*) begin
		main_for_body15_us_us_i_6 = main_entry_coef_out_a;
end
always @(*) begin
	main_for_body15_us_us_i_mul_us_us_i = main_for_body15_us_us_i_mul_us_us_i_stage0_reg;
end
always @(*) begin
		main_for_body15_us_us_i_add23_us_us_i = (main_for_body15_us_us_i_mul_us_us_i + main_for_body15_us_us_i_fir_055_us_us_i_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_12)) begin
		main_for_body15_us_us_i_add23_us_us_i_reg <= main_for_body15_us_us_i_add23_us_us_i;
	end
end
always @(*) begin
		main_for_body15_us_us_i_7 = (main_for_body15_us_us_i_k_154_us_us_i_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_9)) begin
		main_for_body15_us_us_i_7_reg <= main_for_body15_us_us_i_7;
	end
end
always @(*) begin
		main_for_body15_us_us_i_exitcond1 = (main_for_body15_us_us_i_7 == 32'd63);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_9)) begin
		main_for_body15_us_us_i_exitcond1_reg <= main_for_body15_us_us_i_exitcond1;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_inc32_us_i_5) & (fsm_stall == 1'd0)) & (main_for_inc32_us_i_exitcond == 1'd0))) begin
		main_for_cond8_preheader_split_us_us_i_i_058_us_i = main_for_inc32_us_i_1;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_preheader_16) & (fsm_stall == 1'd0))) */ begin
		main_for_cond8_preheader_split_us_us_i_i_058_us_i = 32'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_inc32_us_i_5) & (fsm_stall == 1'd0)) & (main_for_inc32_us_i_exitcond == 1'd0))) begin
		main_for_cond8_preheader_split_us_us_i_i_058_us_i_reg <= main_for_cond8_preheader_split_us_us_i_i_058_us_i;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond8_preheader_split_us_us_i_preheader_16) & (fsm_stall == 1'd0))) begin
		main_for_cond8_preheader_split_us_us_i_i_058_us_i_reg <= main_for_cond8_preheader_split_us_us_i_i_058_us_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_body_i_k_084_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_i_15) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond3_reg == 1'd0))) */ begin
		main_for_body_i_k_084_i = main_for_body_i_8_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_body_i_k_084_i_reg <= main_for_body_i_k_084_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_15) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond3_reg == 1'd0))) begin
		main_for_body_i_k_084_i_reg <= main_for_body_i_k_084_i;
	end
end
always @(*) begin
		main_for_body_i_bit_select = main_for_body_i_k_084_i_reg_width_extended[15:0];
end
always @(*) begin
		main_for_body_i_arrayidx_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_084_i_reg}));
end
always @(*) begin
		main_for_body_i_arrayidx3_i = (1'd0 + (2 * {21'd0,main_for_body_i_k_084_i_reg}));
end
always @(*) begin
		main_for_body_i_8 = ({1'd0,main_for_body_i_k_084_i_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_for_body_i_8_reg <= main_for_body_i_8;
	end
end
always @(*) begin
		main_for_body_i_exitcond3 = (main_for_body_i_8 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_for_body_i_exitcond3_reg <= main_for_body_i_exitcond3;
	end
end
assign main_fir_exit_arrayidx35_i = (1'd0 + (2 * 32'd50));
always @(*) begin
		main_fir_exit_9 = main_entry_vla2_i2_out_a;
end
always @(*) begin
		main_fir_exit_bit_concat = {main_fir_exit_bit_concat_bit_select_operand_0[15:0], main_fir_exit_9[15:0]};
end
always @(*) begin
	main_entry_vla_i1_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_10)) begin
		main_entry_vla_i1_address_a = (main_for_body15_us_us_i_arrayidx17_us_us_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_entry_vla_i1_address_a = (main_for_body_i_arrayidx_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_vla_i1_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_entry_vla_i1_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla_i1_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_entry_vla_i1_in_a = main_for_body_i_bit_select;
	end
end
always @(*) begin
	main_entry_vla2_i2_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_end27_us_us_i_6)) begin
		main_entry_vla2_i2_address_a = (main_for_body15_lr_ph_us_us_i_arrayidx28_us_us_i_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_entry_vla2_i2_address_a = (main_for_body_i_arrayidx3_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_fir_exit_17)) begin
		main_entry_vla2_i2_address_a = (main_fir_exit_arrayidx35_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_vla2_i2_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_end27_us_us_i_6)) begin
		main_entry_vla2_i2_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_entry_vla2_i2_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla2_i2_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_end27_us_us_i_6)) begin
		main_entry_vla2_i2_in_a = main_for_body15_us_us_i_add23_us_us_i_reg;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_14)) begin
		main_entry_vla2_i2_in_a = 16'd0;
	end
end
always @(*) begin
	main_entry_coef_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_coef_address_a = (main_for_body_arrayidx >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body15_us_us_i_10)) begin
		main_entry_coef_address_a = (main_for_body15_us_us_i_arrayidx20_us_us_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_coef_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_coef_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_coef_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_2)) begin
		main_entry_coef_in_a = main_for_body_bit_select1;
	end
end
always @(*) begin
	main_for_body_0_width_extended = {9'd0,main_for_body_0};
end
always @(*) begin
	legup_mult_main_for_body15_us_us_i_mul_us_us_i_en = ~(fsm_stall);
end
always @(posedge clk) begin
	if ((legup_mult_main_for_body15_us_us_i_mul_us_us_i_en == 1'd1)) begin
		main_for_body15_us_us_i_mul_us_us_i_stage0_reg <= (main_for_body15_us_us_i_6 * main_for_body15_us_us_i_5);
	end
end
always @(*) begin
	main_for_body_i_k_084_i_reg_width_extended = {5'd0,main_for_body_i_k_084_i_reg};
end
assign main_fir_exit_bit_concat_bit_select_operand_0 = 16'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_fir_exit_18)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_fir_exit_18)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
