// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Wed Apr 29 09:33:31 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [4:0] LEGUP_0 = 5'd0;
parameter [4:0] LEGUP_F_main_BB_entry_1 = 5'd1;
parameter [4:0] LEGUP_F_main_BB_for_body_i_2 = 5'd2;
parameter [4:0] LEGUP_F_main_BB_for_body_i_3 = 5'd3;
parameter [4:0] LEGUP_F_main_BB_for_body7_i_preheader_4 = 5'd4;
parameter [4:0] LEGUP_F_main_BB_for_body7_i_5 = 5'd5;
parameter [4:0] LEGUP_F_main_BB_for_body7_i_6 = 5'd6;
parameter [4:0] LEGUP_F_main_BB_for_body16_i_preheader_7 = 5'd7;
parameter [4:0] LEGUP_F_main_BB_for_body16_i_8 = 5'd8;
parameter [4:0] LEGUP_F_main_BB_for_body16_i_9 = 5'd9;
parameter [4:0] LEGUP_F_main_BB_for_cond26_preheader_i_preheader_10 = 5'd10;
parameter [4:0] LEGUP_F_main_BB_for_cond26_preheader_i_11 = 5'd11;
parameter [4:0] LEGUP_F_main_BB_for_end59_us_loopexit_i_12 = 5'd12;
parameter [4:0] LEGUP_F_main_BB_for_end59_us_loopexit_i_13 = 5'd13;
parameter [4:0] LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14 = 5'd14;
parameter [4:0] LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15 = 5'd15;
parameter [4:0] LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_16 = 5'd16;
parameter [4:0] LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_17 = 5'd17;
parameter [4:0] LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_18 = 5'd18;
parameter [4:0] LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19 = 5'd19;
parameter [4:0] LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20 = 5'd20;
parameter [4:0] LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_21 = 5'd21;
parameter [4:0] LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_22 = 5'd22;
parameter [4:0] LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_23 = 5'd23;
parameter [4:0] LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24 = 5'd24;
parameter [4:0] LEGUP_F_main_BB_for_inc64_loopexit_i_25 = 5'd25;
parameter [4:0] LEGUP_F_main_BB_kmeans_exit_26 = 5'd26;
parameter [4:0] LEGUP_F_main_BB_kmeans_exit_27 = 5'd27;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [4:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [4:0] next_state;
wire  fsm_stall;
reg [13:0] main_for_body_i_i_0150_i;
reg [13:0] main_for_body_i_i_0150_i_reg;
reg [15:0] main_for_body_i_bit_select11;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx_i;
reg [14:0] main_for_body_i_0;
reg [14:0] main_for_body_i_0_reg;
reg  main_for_body_i_exitcond5;
reg  main_for_body_i_exitcond5_reg;
reg [10:0] main_for_body7_i_i_1148_i;
reg [10:0] main_for_body7_i_i_1148_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body7_i_arrayidx8_i;
reg [11:0] main_for_body7_i_1;
reg [11:0] main_for_body7_i_1_reg;
reg  main_for_body7_i_exitcond;
reg  main_for_body7_i_exitcond_reg;
reg [5:0] main_for_body16_i_i_2147_i;
reg [5:0] main_for_body16_i_i_2147_i_reg;
reg [15:0] main_for_body16_i_bit_select10;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body16_i_arrayidx18_i;
reg [6:0] main_for_body16_i_2;
reg [6:0] main_for_body16_i_2_reg;
reg  main_for_body16_i_exitcond4;
reg  main_for_body16_i_exitcond4_reg;
reg [6:0] main_for_cond26_preheader_i_sp_0145_i;
reg [6:0] main_for_cond26_preheader_i_sp_0145_i_reg;
reg [31:0] main_for_end59_us_loopexit_i_3;
reg [31:0] main_for_end59_us_loopexit_i_3_reg;
reg  main_for_end59_us_loopexit_i_exitcond2;
reg  main_for_end59_us_loopexit_i_exitcond2_reg;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx60_us;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx60_us_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_4;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_4_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var0;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_5;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_5_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var1;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_6;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_6_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var2_reg;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_7;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_7_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var3_reg;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_8;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_8_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var4_reg;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_9;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_9_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var5_reg;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_10;
reg [31:0] main_for_cond35_preheader_lr_ph_us_i_10_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var6_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_pre;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_pre_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_11;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_11_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_12;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_12_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_13;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_13_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_14;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_14_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_15;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_15_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_16;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_16_reg;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_17;
reg [15:0] main_for_cond35_preheader_lr_ph_us_i_17_reg;
reg [31:0] main_for_body38_lr_ph_us_us_i_indvars_iv;
reg [31:0] main_for_body38_lr_ph_us_us_i_indvars_iv_reg;
reg [15:0] main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i;
reg [15:0] main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i_reg;
reg [15:0] main_for_body38_lr_ph_us_us_i_min_0105_us_us_i;
reg [15:0] main_for_body38_lr_ph_us_us_i_min_0105_us_us_i_reg;
reg [15:0] main_for_body38_lr_ph_us_us_i_bit_select9;
reg [15:0] main_for_body38_lr_ph_us_us_i_bit_select9_reg;
reg [28:0] main_for_body38_lr_ph_us_us_i_bit_select;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_1;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_2_reg;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_3_reg;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_4_reg;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_5_reg;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_6_reg;
reg [31:0] main_for_body38_lr_ph_us_us_i_bit_concat1;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_7_reg;
reg [15:0] main_for_body38_lr_ph_us_us_i_18;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i;
reg [15:0] main_for_body38_lr_ph_us_us_i_19;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_1;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i_1;
reg [15:0] main_for_body38_lr_ph_us_us_i_20;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_2;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_2_reg;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i_2;
reg [15:0] main_for_body38_lr_ph_us_us_i_21;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_3;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i_3;
reg [15:0] main_for_body38_lr_ph_us_us_i_22;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_4;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_4_reg;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i_4;
reg [15:0] main_for_body38_lr_ph_us_us_i_23;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_5;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i_5;
reg [15:0] main_for_body38_lr_ph_us_us_i_24;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_6;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_6_reg;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i_6;
reg [15:0] main_for_body38_lr_ph_us_us_i_25;
reg [15:0] main_for_body38_lr_ph_us_us_i_sub_us_us_i_7;
reg [15:0] main_for_body38_lr_ph_us_us_i_add48_us_us_i_7;
reg  main_for_body38_lr_ph_us_us_i_cmp55_us_us_i;
reg [15:0] main_for_body38_lr_ph_us_us_i_min_0_sum_0_us_us_i;
reg [15:0] main_for_body38_lr_ph_us_us_i_min_id_0_c_0_us_us_i;
reg [15:0] main_for_body38_lr_ph_us_us_i_min_id_0_c_0_us_us_i_reg;
reg [31:0] main_for_body38_lr_ph_us_us_i_26;
reg [31:0] main_for_body38_lr_ph_us_us_i_26_reg;
reg  main_for_body38_lr_ph_us_us_i_exitcond1;
reg  main_for_body38_lr_ph_us_us_i_exitcond1_reg;
reg [7:0] main_for_inc64_loopexit_i_27;
reg  main_for_inc64_loopexit_i_exitcond3;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_kmeans_exit_arrayidx67_i;
reg [15:0] main_kmeans_exit_28;
reg [31:0] main_kmeans_exit_bit_concat;
reg [9:0] main_entry_data_out_i_address_a;
reg  main_entry_data_out_i_write_enable_a;
reg [15:0] main_entry_data_out_i_in_a;
wire [15:0] main_entry_data_out_i_out_a;
reg [12:0] main_entry_vla_i1_address_a;
reg  main_entry_vla_i1_write_enable_a;
reg [15:0] main_entry_vla_i1_in_a;
wire [15:0] main_entry_vla_i1_out_a;
reg [12:0] main_entry_vla_i1_address_b;
wire  main_entry_vla_i1_write_enable_b;
wire [15:0] main_entry_vla_i1_in_b;
wire [15:0] main_entry_vla_i1_out_b;
reg [5:0] main_entry_vla2_i2_address_a;
reg  main_entry_vla2_i2_write_enable_a;
reg [15:0] main_entry_vla2_i2_in_a;
wire [15:0] main_entry_vla2_i2_out_a;
reg [5:0] main_entry_vla2_i2_address_b;
wire  main_entry_vla2_i2_write_enable_b;
wire [15:0] main_entry_vla2_i2_in_b;
wire [15:0] main_entry_vla2_i2_out_b;
reg [15:0] main_for_body_i_i_0150_i_reg_width_extended;
reg [15:0] main_for_body16_i_i_2147_i_reg_width_extended;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat8_bit_select_operand_2;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat7_bit_select_operand_2;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat6_bit_select_operand_2;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat5_bit_select_operand_2;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat4_bit_select_operand_2;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat3_bit_select_operand_2;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat2_bit_select_operand_2;
wire [2:0] main_for_body38_lr_ph_us_us_i_bit_concat1_bit_select_operand_2;
wire [15:0] main_kmeans_exit_bit_concat_bit_select_operand_0;



//   %data_out.i = alloca [1024 x i16], align 2, !dbg !46, !MSB !47, !LSB !48, !extendFrom !47
ram_single_port main_entry_data_out_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_data_out_i_address_a ),
	.wren_a( main_entry_data_out_i_write_enable_a ),
	.data_a( main_entry_data_out_i_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_data_out_i_out_a )
);
defparam main_entry_data_out_i.width_a = 16;
defparam main_entry_data_out_i.widthad_a = 10;
defparam main_entry_data_out_i.width_be_a = 2;
defparam main_entry_data_out_i.numwords_a = 1024;
defparam main_entry_data_out_i.latency = 1;


//   %vla.i1 = alloca [8192 x i16], align 2, !dbg !49, !MSB !47, !LSB !48, !extendFrom !47
ram_dual_port main_entry_vla_i1 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla_i1_address_a ),
	.wren_a( main_entry_vla_i1_write_enable_a ),
	.data_a( main_entry_vla_i1_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_vla_i1_out_a ),
	.address_b( main_entry_vla_i1_address_b ),
	.wren_b( main_entry_vla_i1_write_enable_b ),
	.data_b( main_entry_vla_i1_in_b ),
	.byteena_b( {2{1'b1}} ),
	.q_b( main_entry_vla_i1_out_b )
);
defparam main_entry_vla_i1.width_a = 16;
defparam main_entry_vla_i1.widthad_a = 13;
defparam main_entry_vla_i1.width_be_a = 2;
defparam main_entry_vla_i1.numwords_a = 8192;
defparam main_entry_vla_i1.width_b = 16;
defparam main_entry_vla_i1.widthad_b = 13;
defparam main_entry_vla_i1.width_be_b = 2;
defparam main_entry_vla_i1.numwords_b = 8192;
defparam main_entry_vla_i1.latency = 1;


//   %vla2.i2 = alloca [40 x i16], align 2, !dbg !50, !MSB !47, !LSB !48, !extendFrom !47
ram_dual_port main_entry_vla2_i2 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla2_i2_address_a ),
	.wren_a( main_entry_vla2_i2_write_enable_a ),
	.data_a( main_entry_vla2_i2_in_a ),
	.byteena_a( {2{1'b1}} ),
	.q_a( main_entry_vla2_i2_out_a ),
	.address_b( main_entry_vla2_i2_address_b ),
	.wren_b( main_entry_vla2_i2_write_enable_b ),
	.data_b( main_entry_vla2_i2_in_b ),
	.byteena_b( {2{1'b1}} ),
	.q_b( main_entry_vla2_i2_out_b )
);
defparam main_entry_vla2_i2.width_a = 16;
defparam main_entry_vla2_i2.widthad_a = 6;
defparam main_entry_vla2_i2.width_be_a = 2;
defparam main_entry_vla2_i2.numwords_a = 40;
defparam main_entry_vla2_i2.width_b = 16;
defparam main_entry_vla2_i2.widthad_b = 6;
defparam main_entry_vla2_i2.width_be_b = 2;
defparam main_entry_vla2_i2.numwords_b = 40;
defparam main_entry_vla2_i2.latency = 1;

/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_kmeans_exit_27)) begin
		$write("%d\n", $signed(main_kmeans_exit_bit_concat));
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_for_body_i_2;
LEGUP_F_main_BB_for_body16_i_8:
		next_state = LEGUP_F_main_BB_for_body16_i_9;
LEGUP_F_main_BB_for_body16_i_9:
	if ((fsm_stall == 1'd0) && (main_for_body16_i_exitcond4_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond26_preheader_i_preheader_10;
	else if ((fsm_stall == 1'd0) && (main_for_body16_i_exitcond4_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body16_i_8;
LEGUP_F_main_BB_for_body16_i_preheader_7:
		next_state = LEGUP_F_main_BB_for_body16_i_8;
LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20:
		next_state = LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_21;
LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_21:
		next_state = LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_22;
LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_22:
		next_state = LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_23;
LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_23:
		next_state = LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24;
LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24:
	if ((fsm_stall == 1'd0) && (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_end59_us_loopexit_i_12;
	else if ((fsm_stall == 1'd0) && (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20;
LEGUP_F_main_BB_for_body7_i_5:
		next_state = LEGUP_F_main_BB_for_body7_i_6;
LEGUP_F_main_BB_for_body7_i_6:
	if ((fsm_stall == 1'd0) && (main_for_body7_i_exitcond_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_body16_i_preheader_7;
	else if ((fsm_stall == 1'd0) && (main_for_body7_i_exitcond_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body7_i_5;
LEGUP_F_main_BB_for_body7_i_preheader_4:
		next_state = LEGUP_F_main_BB_for_body7_i_5;
LEGUP_F_main_BB_for_body_i_2:
		next_state = LEGUP_F_main_BB_for_body_i_3;
LEGUP_F_main_BB_for_body_i_3:
	if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond5_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_body7_i_preheader_4;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond5_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_2;
LEGUP_F_main_BB_for_cond26_preheader_i_11:
		next_state = LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14;
LEGUP_F_main_BB_for_cond26_preheader_i_preheader_10:
		next_state = LEGUP_F_main_BB_for_cond26_preheader_i_11;
LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14:
		next_state = LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15;
LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15:
		next_state = LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_16;
LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_16:
		next_state = LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_17;
LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_17:
		next_state = LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_18;
LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_18:
		next_state = LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19;
LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19:
		next_state = LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20;
LEGUP_F_main_BB_for_end59_us_loopexit_i_12:
		next_state = LEGUP_F_main_BB_for_end59_us_loopexit_i_13;
LEGUP_F_main_BB_for_end59_us_loopexit_i_13:
	if ((fsm_stall == 1'd0) && (main_for_end59_us_loopexit_i_exitcond2_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc64_loopexit_i_25;
	else if ((fsm_stall == 1'd0) && (main_for_end59_us_loopexit_i_exitcond2_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14;
LEGUP_F_main_BB_for_inc64_loopexit_i_25:
	if ((fsm_stall == 1'd0) && (main_for_inc64_loopexit_i_exitcond3 == 1'd1))
		next_state = LEGUP_F_main_BB_kmeans_exit_26;
	else if ((fsm_stall == 1'd0) && (main_for_inc64_loopexit_i_exitcond3 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond26_preheader_i_11;
LEGUP_F_main_BB_kmeans_exit_26:
		next_state = LEGUP_F_main_BB_kmeans_exit_27;
LEGUP_F_main_BB_kmeans_exit_27:
		next_state = LEGUP_0;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_0150_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_i_3) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond5_reg == 1'd0))) */ begin
		main_for_body_i_i_0150_i = main_for_body_i_0_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_0150_i_reg <= main_for_body_i_i_0150_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_3) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond5_reg == 1'd0))) begin
		main_for_body_i_i_0150_i_reg <= main_for_body_i_i_0150_i;
	end
end
always @(*) begin
		main_for_body_i_bit_select11 = main_for_body_i_i_0150_i_reg_width_extended[15:0];
end
always @(*) begin
		main_for_body_i_arrayidx_i = (1'd0 + (2 * {18'd0,main_for_body_i_i_0150_i_reg}));
end
always @(*) begin
		main_for_body_i_0 = ({1'd0,main_for_body_i_i_0150_i_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_for_body_i_0_reg <= main_for_body_i_0;
	end
end
always @(*) begin
		main_for_body_i_exitcond5 = (main_for_body_i_0 == 32'd8192);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_for_body_i_exitcond5_reg <= main_for_body_i_exitcond5;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body7_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_body7_i_i_1148_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body7_i_6) & (fsm_stall == 1'd0)) & (main_for_body7_i_exitcond_reg == 1'd0))) */ begin
		main_for_body7_i_i_1148_i = main_for_body7_i_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body7_i_preheader_4) & (fsm_stall == 1'd0))) begin
		main_for_body7_i_i_1148_i_reg <= main_for_body7_i_i_1148_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body7_i_6) & (fsm_stall == 1'd0)) & (main_for_body7_i_exitcond_reg == 1'd0))) begin
		main_for_body7_i_i_1148_i_reg <= main_for_body7_i_i_1148_i;
	end
end
always @(*) begin
		main_for_body7_i_arrayidx8_i = (1'd0 + (2 * {21'd0,main_for_body7_i_i_1148_i_reg}));
end
always @(*) begin
		main_for_body7_i_1 = ({1'd0,main_for_body7_i_i_1148_i_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body7_i_5)) begin
		main_for_body7_i_1_reg <= main_for_body7_i_1;
	end
end
always @(*) begin
		main_for_body7_i_exitcond = (main_for_body7_i_1 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body7_i_5)) begin
		main_for_body7_i_exitcond_reg <= main_for_body7_i_exitcond;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body16_i_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_body16_i_i_2147_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body16_i_9) & (fsm_stall == 1'd0)) & (main_for_body16_i_exitcond4_reg == 1'd0))) */ begin
		main_for_body16_i_i_2147_i = main_for_body16_i_2_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body16_i_preheader_7) & (fsm_stall == 1'd0))) begin
		main_for_body16_i_i_2147_i_reg <= main_for_body16_i_i_2147_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body16_i_9) & (fsm_stall == 1'd0)) & (main_for_body16_i_exitcond4_reg == 1'd0))) begin
		main_for_body16_i_i_2147_i_reg <= main_for_body16_i_i_2147_i;
	end
end
always @(*) begin
		main_for_body16_i_bit_select10 = main_for_body16_i_i_2147_i_reg_width_extended[15:0];
end
always @(*) begin
		main_for_body16_i_arrayidx18_i = (1'd0 + (2 * {26'd0,main_for_body16_i_i_2147_i_reg}));
end
always @(*) begin
		main_for_body16_i_2 = ({1'd0,main_for_body16_i_i_2147_i_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body16_i_8)) begin
		main_for_body16_i_2_reg <= main_for_body16_i_2;
	end
end
always @(*) begin
		main_for_body16_i_exitcond4 = (main_for_body16_i_2 == 32'd40);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body16_i_8)) begin
		main_for_body16_i_exitcond4_reg <= main_for_body16_i_exitcond4;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond26_preheader_i_preheader_10) & (fsm_stall == 1'd0))) begin
		main_for_cond26_preheader_i_sp_0145_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc64_loopexit_i_25) & (fsm_stall == 1'd0)) & (main_for_inc64_loopexit_i_exitcond3 == 1'd0))) */ begin
		main_for_cond26_preheader_i_sp_0145_i = main_for_inc64_loopexit_i_27;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond26_preheader_i_preheader_10) & (fsm_stall == 1'd0))) begin
		main_for_cond26_preheader_i_sp_0145_i_reg <= main_for_cond26_preheader_i_sp_0145_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc64_loopexit_i_25) & (fsm_stall == 1'd0)) & (main_for_inc64_loopexit_i_exitcond3 == 1'd0))) begin
		main_for_cond26_preheader_i_sp_0145_i_reg <= main_for_cond26_preheader_i_sp_0145_i;
	end
end
always @(*) begin
		main_for_end59_us_loopexit_i_3 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_end59_us_loopexit_i_12)) begin
		main_for_end59_us_loopexit_i_3_reg <= main_for_end59_us_loopexit_i_3;
	end
end
always @(*) begin
		main_for_end59_us_loopexit_i_exitcond2 = (main_for_end59_us_loopexit_i_3 == 32'd1024);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_end59_us_loopexit_i_12)) begin
		main_for_end59_us_loopexit_i_exitcond2_reg <= main_for_end59_us_loopexit_i_exitcond2;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond26_preheader_i_11) & (fsm_stall == 1'd0))) begin
		main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_end59_us_loopexit_i_13) & (fsm_stall == 1'd0)) & (main_for_end59_us_loopexit_i_exitcond2_reg == 1'd0))) */ begin
		main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i = main_for_end59_us_loopexit_i_3_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond26_preheader_i_11) & (fsm_stall == 1'd0))) begin
		main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg <= main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_end59_us_loopexit_i_13) & (fsm_stall == 1'd0)) & (main_for_end59_us_loopexit_i_exitcond2_reg == 1'd0))) begin
		main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg <= main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx60_us = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx60_us_reg <= main_for_cond35_preheader_lr_ph_us_i_arrayidx60_us;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg));
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_4 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd8);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_4_reg <= main_for_cond35_preheader_lr_ph_us_i_4;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var0 = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_4_reg));
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_5 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd16);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_5_reg <= main_for_cond35_preheader_lr_ph_us_i_5;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var1 = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_5_reg));
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_6 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd24);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_6_reg <= main_for_cond35_preheader_lr_ph_us_i_6;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var2 = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_6_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var2_reg <= main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var2;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_7 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd32);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_7_reg <= main_for_cond35_preheader_lr_ph_us_i_7;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var3 = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_7_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var3_reg <= main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var3;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_8 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd40);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_8_reg <= main_for_cond35_preheader_lr_ph_us_i_8;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var4 = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_8_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var4_reg <= main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var4;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_9 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd48);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_9_reg <= main_for_cond35_preheader_lr_ph_us_i_9;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var5 = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_9_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var5_reg <= main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var5;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_10 = (main_for_cond35_preheader_lr_ph_us_i_i_3109_us_i_reg + 32'd56);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_for_cond35_preheader_lr_ph_us_i_10_reg <= main_for_cond35_preheader_lr_ph_us_i_10;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var6 = (1'd0 + (2 * main_for_cond35_preheader_lr_ph_us_i_10_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var6_reg <= main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var6;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_pre = main_entry_vla_i1_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_for_cond35_preheader_lr_ph_us_i_pre_reg <= main_for_cond35_preheader_lr_ph_us_i_pre;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_11 = main_entry_vla_i1_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_16)) begin
		main_for_cond35_preheader_lr_ph_us_i_11_reg <= main_for_cond35_preheader_lr_ph_us_i_11;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_12 = main_entry_vla_i1_out_b;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_16)) begin
		main_for_cond35_preheader_lr_ph_us_i_12_reg <= main_for_cond35_preheader_lr_ph_us_i_12;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_13 = main_entry_vla_i1_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_17)) begin
		main_for_cond35_preheader_lr_ph_us_i_13_reg <= main_for_cond35_preheader_lr_ph_us_i_13;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_14 = main_entry_vla_i1_out_b;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_17)) begin
		main_for_cond35_preheader_lr_ph_us_i_14_reg <= main_for_cond35_preheader_lr_ph_us_i_14;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_15 = main_entry_vla_i1_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_18)) begin
		main_for_cond35_preheader_lr_ph_us_i_15_reg <= main_for_cond35_preheader_lr_ph_us_i_15;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_16 = main_entry_vla_i1_out_b;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_18)) begin
		main_for_cond35_preheader_lr_ph_us_i_16_reg <= main_for_cond35_preheader_lr_ph_us_i_16;
	end
end
always @(*) begin
		main_for_cond35_preheader_lr_ph_us_i_17 = main_entry_vla_i1_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19)) begin
		main_for_cond35_preheader_lr_ph_us_i_17_reg <= main_for_cond35_preheader_lr_ph_us_i_17;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19) & (fsm_stall == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_indvars_iv = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24) & (fsm_stall == 1'd0)) & (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd0))) */ begin
		main_for_body38_lr_ph_us_us_i_indvars_iv = main_for_body38_lr_ph_us_us_i_26_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19) & (fsm_stall == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_indvars_iv_reg <= main_for_body38_lr_ph_us_us_i_indvars_iv;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24) & (fsm_stall == 1'd0)) & (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_indvars_iv_reg <= main_for_body38_lr_ph_us_us_i_indvars_iv;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19) & (fsm_stall == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i = 16'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24) & (fsm_stall == 1'd0)) & (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd0))) */ begin
		main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i = main_for_body38_lr_ph_us_us_i_min_id_0_c_0_us_us_i;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19) & (fsm_stall == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i_reg <= main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24) & (fsm_stall == 1'd0)) & (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i_reg <= main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19) & (fsm_stall == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_min_0105_us_us_i = -16'd32203;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24) & (fsm_stall == 1'd0)) & (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd0))) */ begin
		main_for_body38_lr_ph_us_us_i_min_0105_us_us_i = main_for_body38_lr_ph_us_us_i_min_0_sum_0_us_us_i;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_19) & (fsm_stall == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_min_0105_us_us_i_reg <= main_for_body38_lr_ph_us_us_i_min_0105_us_us_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24) & (fsm_stall == 1'd0)) & (main_for_body38_lr_ph_us_us_i_exitcond1_reg == 1'd0))) begin
		main_for_body38_lr_ph_us_us_i_min_0105_us_us_i_reg <= main_for_body38_lr_ph_us_us_i_min_0105_us_us_i;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_select9 = main_for_body38_lr_ph_us_us_i_indvars_iv_reg[15:0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_bit_select9_reg <= main_for_body38_lr_ph_us_us_i_bit_select9;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_select = main_for_body38_lr_ph_us_us_i_indvars_iv_reg[28:0];
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat8 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat8_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat8));
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat7 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat7_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_1 = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat7));
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat6 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat6_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_2 = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat6));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_2_reg <= main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_2;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat5 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat5_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_3 = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat5));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_3_reg <= main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_3;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat4 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat4_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_4 = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat4));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_4_reg <= main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_4;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat3 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat3_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_5 = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat3));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_5_reg <= main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_5;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat2 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat2_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_6 = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat2));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_6_reg <= main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_6;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_bit_concat1 = {main_for_body38_lr_ph_us_us_i_bit_select[28:0], main_for_body38_lr_ph_us_us_i_bit_concat1_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_7 = (1'd0 + (2 * main_for_body38_lr_ph_us_us_i_bit_concat1));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_7_reg <= main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_7;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_18 = main_entry_vla2_i2_out_a;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i = (main_for_cond35_preheader_lr_ph_us_i_pre_reg - main_for_body38_lr_ph_us_us_i_18);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_19 = main_entry_vla2_i2_out_b;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_1 = (main_for_cond35_preheader_lr_ph_us_i_11_reg + main_for_body38_lr_ph_us_us_i_add48_us_us_i);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i_1 = (main_for_body38_lr_ph_us_us_i_sub_us_us_i_1 - main_for_body38_lr_ph_us_us_i_19);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_20 = main_entry_vla2_i2_out_a;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_2 = (main_for_cond35_preheader_lr_ph_us_i_12_reg + main_for_body38_lr_ph_us_us_i_add48_us_us_i_1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_21)) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_2_reg <= main_for_body38_lr_ph_us_us_i_sub_us_us_i_2;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i_2 = (main_for_body38_lr_ph_us_us_i_sub_us_us_i_2_reg - main_for_body38_lr_ph_us_us_i_20);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_21 = main_entry_vla2_i2_out_b;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_3 = (main_for_cond35_preheader_lr_ph_us_i_13_reg + main_for_body38_lr_ph_us_us_i_add48_us_us_i_2);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i_3 = (main_for_body38_lr_ph_us_us_i_sub_us_us_i_3 - main_for_body38_lr_ph_us_us_i_21);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_22 = main_entry_vla2_i2_out_a;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_4 = (main_for_cond35_preheader_lr_ph_us_i_14_reg + main_for_body38_lr_ph_us_us_i_add48_us_us_i_3);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_22)) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_4_reg <= main_for_body38_lr_ph_us_us_i_sub_us_us_i_4;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i_4 = (main_for_body38_lr_ph_us_us_i_sub_us_us_i_4_reg - main_for_body38_lr_ph_us_us_i_22);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_23 = main_entry_vla2_i2_out_b;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_5 = (main_for_cond35_preheader_lr_ph_us_i_15_reg + main_for_body38_lr_ph_us_us_i_add48_us_us_i_4);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i_5 = (main_for_body38_lr_ph_us_us_i_sub_us_us_i_5 - main_for_body38_lr_ph_us_us_i_23);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_24 = main_entry_vla2_i2_out_a;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_6 = (main_for_cond35_preheader_lr_ph_us_i_16_reg + main_for_body38_lr_ph_us_us_i_add48_us_us_i_5);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_23)) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_6_reg <= main_for_body38_lr_ph_us_us_i_sub_us_us_i_6;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i_6 = (main_for_body38_lr_ph_us_us_i_sub_us_us_i_6_reg - main_for_body38_lr_ph_us_us_i_24);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_25 = main_entry_vla2_i2_out_b;
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_sub_us_us_i_7 = (main_for_cond35_preheader_lr_ph_us_i_17_reg + main_for_body38_lr_ph_us_us_i_add48_us_us_i_6);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_add48_us_us_i_7 = (main_for_body38_lr_ph_us_us_i_sub_us_us_i_7 - main_for_body38_lr_ph_us_us_i_25);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_cmp55_us_us_i = (main_for_body38_lr_ph_us_us_i_add48_us_us_i_7 > main_for_body38_lr_ph_us_us_i_min_0105_us_us_i_reg);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_min_0_sum_0_us_us_i = (main_for_body38_lr_ph_us_us_i_cmp55_us_us_i ? main_for_body38_lr_ph_us_us_i_min_0105_us_us_i_reg : main_for_body38_lr_ph_us_us_i_add48_us_us_i_7);
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_min_id_0_c_0_us_us_i = (main_for_body38_lr_ph_us_us_i_cmp55_us_us_i ? main_for_body38_lr_ph_us_us_i_min_id_0106_us_us_i_reg : main_for_body38_lr_ph_us_us_i_bit_select9_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_24)) begin
		main_for_body38_lr_ph_us_us_i_min_id_0_c_0_us_us_i_reg <= main_for_body38_lr_ph_us_us_i_min_id_0_c_0_us_us_i;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_26 = (main_for_body38_lr_ph_us_us_i_indvars_iv_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_26_reg <= main_for_body38_lr_ph_us_us_i_26;
	end
end
always @(*) begin
		main_for_body38_lr_ph_us_us_i_exitcond1 = (main_for_body38_lr_ph_us_us_i_26 == 32'd5);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_for_body38_lr_ph_us_us_i_exitcond1_reg <= main_for_body38_lr_ph_us_us_i_exitcond1;
	end
end
always @(*) begin
		main_for_inc64_loopexit_i_27 = ({1'd0,main_for_cond26_preheader_i_sp_0145_i_reg} + 32'd1);
end
always @(*) begin
		main_for_inc64_loopexit_i_exitcond3 = (main_for_inc64_loopexit_i_27 == 32'd100);
end
assign main_kmeans_exit_arrayidx67_i = (1'd0 + (2 * 32'd50));
always @(*) begin
		main_kmeans_exit_28 = main_entry_data_out_i_out_a;
end
always @(*) begin
		main_kmeans_exit_bit_concat = {main_kmeans_exit_bit_concat_bit_select_operand_0[15:0], main_kmeans_exit_28[15:0]};
end
always @(*) begin
	main_entry_data_out_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body7_i_5)) begin
		main_entry_data_out_i_address_a = (main_for_body7_i_arrayidx8_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_end59_us_loopexit_i_12)) begin
		main_entry_data_out_i_address_a = (main_for_cond35_preheader_lr_ph_us_i_arrayidx60_us_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_kmeans_exit_26)) begin
		main_entry_data_out_i_address_a = (main_kmeans_exit_arrayidx67_i >>> 3'd1);
	end
end
always @(*) begin
	main_entry_data_out_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body7_i_5)) begin
		main_entry_data_out_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end59_us_loopexit_i_12)) begin
		main_entry_data_out_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_data_out_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body7_i_5)) begin
		main_entry_data_out_i_in_a = 16'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end59_us_loopexit_i_12)) begin
		main_entry_data_out_i_in_a = main_for_body38_lr_ph_us_us_i_min_id_0_c_0_us_us_i_reg;
	end
end
always @(*) begin
	main_entry_vla_i1_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_vla_i1_address_a = (main_for_body_i_arrayidx_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_14)) begin
		main_entry_vla_i1_address_a = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_entry_vla_i1_address_a = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var0 >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_16)) begin
		main_entry_vla_i1_address_a = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var2_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_17)) begin
		main_entry_vla_i1_address_a = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var4_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_18)) begin
		main_entry_vla_i1_address_a = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var6_reg >>> 3'd1);
	end
end
always @(*) begin
	main_entry_vla_i1_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_vla_i1_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla_i1_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_2)) begin
		main_entry_vla_i1_in_a = main_for_body_i_bit_select11;
	end
end
always @(*) begin
	main_entry_vla_i1_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_15)) begin
		main_entry_vla_i1_address_b = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var1 >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_16)) begin
		main_entry_vla_i1_address_b = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var3_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond35_preheader_lr_ph_us_i_17)) begin
		main_entry_vla_i1_address_b = (main_for_cond35_preheader_lr_ph_us_i_arrayidx40_us_var5_reg >>> 3'd1);
	end
end
assign main_entry_vla_i1_write_enable_b = 'd0;
assign main_entry_vla_i1_in_b = 'dx;
always @(*) begin
	main_entry_vla2_i2_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body16_i_8)) begin
		main_entry_vla2_i2_address_a = (main_for_body16_i_arrayidx18_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_entry_vla2_i2_address_a = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_21)) begin
		main_entry_vla2_i2_address_a = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_2_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_22)) begin
		main_entry_vla2_i2_address_a = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_4_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_23)) begin
		main_entry_vla2_i2_address_a = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_6_reg >>> 3'd1);
	end
end
always @(*) begin
	main_entry_vla2_i2_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body16_i_8)) begin
		main_entry_vla2_i2_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla2_i2_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body16_i_8)) begin
		main_entry_vla2_i2_in_a = main_for_body16_i_bit_select10;
	end
end
always @(*) begin
	main_entry_vla2_i2_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_20)) begin
		main_entry_vla2_i2_address_b = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_1 >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_21)) begin
		main_entry_vla2_i2_address_b = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_3_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_22)) begin
		main_entry_vla2_i2_address_b = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_5_reg >>> 3'd1);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body38_lr_ph_us_us_i_23)) begin
		main_entry_vla2_i2_address_b = (main_for_body38_lr_ph_us_us_i_arrayidx45_us_us_i_7_reg >>> 3'd1);
	end
end
assign main_entry_vla2_i2_write_enable_b = 'd0;
assign main_entry_vla2_i2_in_b = 'dx;
always @(*) begin
	main_for_body_i_i_0150_i_reg_width_extended = {2'd0,main_for_body_i_i_0150_i_reg};
end
always @(*) begin
	main_for_body16_i_i_2147_i_reg_width_extended = {10'd0,main_for_body16_i_i_2147_i_reg};
end
assign main_for_body38_lr_ph_us_us_i_bit_concat8_bit_select_operand_2 = 3'd0;
assign main_for_body38_lr_ph_us_us_i_bit_concat7_bit_select_operand_2 = 3'd1;
assign main_for_body38_lr_ph_us_us_i_bit_concat6_bit_select_operand_2 = 3'd2;
assign main_for_body38_lr_ph_us_us_i_bit_concat5_bit_select_operand_2 = 3'd3;
assign main_for_body38_lr_ph_us_us_i_bit_concat4_bit_select_operand_2 = -3'd4;
assign main_for_body38_lr_ph_us_us_i_bit_concat3_bit_select_operand_2 = -3'd3;
assign main_for_body38_lr_ph_us_us_i_bit_concat2_bit_select_operand_2 = -3'd2;
assign main_for_body38_lr_ph_us_us_i_bit_concat1_bit_select_operand_2 = -3'd1;
assign main_kmeans_exit_bit_concat_bit_select_operand_0 = 16'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_kmeans_exit_27)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_kmeans_exit_27)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a,
	address_b,
	wren_b,
	data_b,
	byteena_b,
	q_b
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_be_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  width_be_b = 1'd0;
parameter  init_file_mem = {`MEM_INIT_DIR, "UNUSED.mem"};
parameter  latency = 1;

input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
reg [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
reg [(width_b-1):0] q_b_wire;
input  wren_b;
input [(width_a-1):0] data_b;
input [width_be_a-1:0] byteena_b;

reg [width_a-1:0] ram [numwords_a-1:0];

initial begin
	if (init_file_mem != {`MEM_INIT_DIR, "UNUSED.mem"})
        $readmemb(init_file_mem, ram);
end

localparam input_latency = ((latency - 1) >> 1);
localparam output_latency = (latency - 1) - input_latency;
integer j;

reg [(widthad_a-1):0] address_a_reg[input_latency:0];
reg  wren_a_reg[input_latency:0];
reg [(width_a-1):0] data_a_reg[input_latency:0];
reg [(width_be_a-1):0] byteena_a_reg[input_latency:0];
reg [(widthad_b-1):0] address_b_reg[input_latency:0];
reg  wren_b_reg[input_latency:0];
reg [(width_b-1):0] data_b_reg[input_latency:0];
reg [(width_be_b-1):0] byteena_b_reg[input_latency:0];

always @(*)
begin
  address_a_reg[0] = address_a;
  wren_a_reg[0] = wren_a;
  data_a_reg[0] = data_a;
  byteena_a_reg[0] = byteena_a;
  address_b_reg[0] = address_b;
  wren_b_reg[0] = wren_b;
  data_b_reg[0] = data_b;
  byteena_b_reg[0] = byteena_b;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < input_latency; j=j+1)
   begin
       address_a_reg[j+1] <= address_a_reg[j];
       wren_a_reg[j+1] <= wren_a_reg[j];
       data_a_reg[j+1] <= data_a_reg[j];
       byteena_a_reg[j+1] <= byteena_a_reg[j];
       address_b_reg[j+1] <= address_b_reg[j];
       wren_b_reg[j+1] <= wren_b_reg[j];
       data_b_reg[j+1] <= data_b_reg[j];
       byteena_b_reg[j+1] <= byteena_b_reg[j];
   end
end

always @ (posedge clk)
begin
    if (clken)
    begin // Port a
        if (wren_a_reg[input_latency])
        begin
            ram[address_a_reg[input_latency]] <= data_a_reg[input_latency];
            q_a_wire <= data_a_reg[input_latency];
        end
        else begin
            q_a_wire <= ram[address_a_reg[input_latency]];
        end
    end
end

always @ (posedge clk)
begin
    if (clken)
    begin // Port b
        if (wren_b_reg[input_latency])
        begin
            ram[address_b_reg[input_latency]] <= data_b_reg[input_latency];
            q_b_wire <= data_b_reg[input_latency];
        end
        else begin
            q_b_wire <= ram[address_b_reg[input_latency]];
        end
    end
end


reg [(width_a-1):0] q_a_reg[output_latency:0];

always @(*)
begin
   q_a_reg[0] <= q_a_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_a_reg[j+1] <= q_a_reg[j];
   end
end

assign q_a = q_a_reg[output_latency];
reg [(width_b-1):0] q_b_reg[output_latency:0];

always @(*)
begin
   q_b_reg[0] <= q_b_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_b_reg[j+1] <= q_b_reg[j];
   end
end

assign q_b = q_b_reg[output_latency];

endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
