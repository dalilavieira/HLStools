// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Mon May  4 13:14:12 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [3:0] LEGUP_0 = 4'd0;
parameter [3:0] LEGUP_F_main_BB_while_body_lr_ph_i_1 = 4'd1;
parameter [3:0] LEGUP_F_main_BB_while_cond_i_2 = 4'd2;
parameter [3:0] LEGUP_F_main_BB_while_body_i_3 = 4'd3;
parameter [3:0] LEGUP_F_main_BB_while_body_i_4 = 4'd4;
parameter [3:0] LEGUP_F_main_BB_if_else_i_5 = 4'd5;
parameter [3:0] LEGUP_F_main_BB_mmc_exit_loopexit_6 = 4'd6;
parameter [3:0] LEGUP_F_main_BB_mmc_exit_loopexit1_7 = 4'd7;
parameter [3:0] LEGUP_F_main_BB_mmc_exit_8 = 4'd8;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [3:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [3:0] next_state;
wire  fsm_stall;
reg [31:0] main_while_body_lr_ph_i_indvar3;
reg [31:0] main_while_body_lr_ph_i_indvar3_reg;
reg [31:0] main_while_body_lr_ph_i_F2_0_ph15_i;
reg [31:0] main_while_body_lr_ph_i_F2_0_ph15_i_reg;
reg [30:0] main_while_body_lr_ph_i_bit_select3;
reg [29:0] main_while_body_lr_ph_i_bit_select1;
reg [31:0] main_while_body_lr_ph_i_bit_concat4;
reg [31:0] main_while_body_lr_ph_i_bit_concat2;
reg [31:0] main_while_body_lr_ph_i_sr_add;
reg [31:0] main_while_body_lr_ph_i_add2_i;
reg [31:0] main_while_body_lr_ph_i_add2_i_reg;
reg [31:0] main_while_body_lr_ph_i_F1_0_ph14_i;
reg [31:0] main_while_body_lr_ph_i_F1_0_ph14_i_reg;
reg [31:0] main_while_body_lr_ph_i_0;
reg [31:0] main_while_body_lr_ph_i_0_reg;
reg [31:0] main_while_cond_i_add_i;
reg  main_while_cond_i_cmp_i;
reg [31:0] main_while_cond_i_indvar_next;
reg [31:0] main_while_body_i_indvar;
reg [31:0] main_while_body_i_indvar_reg;
reg [28:0] main_while_body_i_bit_select;
reg [31:0] main_while_body_i_sr_negate;
reg [31:0] main_while_body_i_bit_concat;
reg [31:0] main_while_body_i_sr_add7;
reg [31:0] main_while_body_i_sr_add7_reg;
reg [31:0] main_while_body_i_F2_011_i;
reg [31:0] main_while_body_i_F2_011_i_reg;
reg  main_while_body_i_cmp1_i;
reg  main_if_else_i_cmp10_i;
reg [31:0] main_if_else_i_indvar_next4;
reg [31:0] main_mmc_exit_F1_0_ph_lcssa_i;
reg [31:0] main_mmc_exit_F1_0_ph_lcssa_i_reg;
wire  main_while_body_lr_ph_i_bit_concat4_bit_select_operand_2;
wire [1:0] main_while_body_lr_ph_i_bit_concat2_bit_select_operand_2;
wire [2:0] main_while_body_i_bit_concat_bit_select_operand_2;


/* Unsynthesizable Statements */
/* synthesis translate_off */
always @(posedge clk)
	if (!fsm_stall) begin
	if ((cur_state == LEGUP_F_main_BB_mmc_exit_8)) begin
		$write("mmc of %d and %d is %d\n", 32'd6, 32'd7, $signed(main_mmc_exit_F1_0_ph_lcssa_i_reg));
		// to fix quartus warning
		if (reset == 1'b0 && ^(32'd6) === 1'bX) finish <= 0;
		if (reset == 1'b0 && ^(32'd7) === 1'bX) finish <= 0;
		if (reset == 1'b0 && ^(main_mmc_exit_F1_0_ph_lcssa_i_reg) === 1'bX) finish <= 0;
	end
end
/* synthesis translate_on */
always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_while_body_lr_ph_i_1;
LEGUP_F_main_BB_if_else_i_5:
	if ((fsm_stall == 1'd0) && (main_if_else_i_cmp10_i == 1'd1))
		next_state = LEGUP_F_main_BB_mmc_exit_loopexit1_7;
	else if ((fsm_stall == 1'd0) && (main_if_else_i_cmp10_i == 1'd0))
		next_state = LEGUP_F_main_BB_while_body_lr_ph_i_1;
LEGUP_F_main_BB_mmc_exit_8:
		next_state = LEGUP_0;
LEGUP_F_main_BB_mmc_exit_loopexit1_7:
		next_state = LEGUP_F_main_BB_mmc_exit_8;
LEGUP_F_main_BB_mmc_exit_loopexit_6:
		next_state = LEGUP_F_main_BB_mmc_exit_8;
LEGUP_F_main_BB_while_body_i_3:
		next_state = LEGUP_F_main_BB_while_body_i_4;
LEGUP_F_main_BB_while_body_i_4:
	if ((fsm_stall == 1'd0) && (main_while_body_i_cmp1_i == 1'd1))
		next_state = LEGUP_F_main_BB_while_cond_i_2;
	else if ((fsm_stall == 1'd0) && (main_while_body_i_cmp1_i == 1'd0))
		next_state = LEGUP_F_main_BB_if_else_i_5;
LEGUP_F_main_BB_while_body_lr_ph_i_1:
		next_state = LEGUP_F_main_BB_while_body_i_3;
LEGUP_F_main_BB_while_cond_i_2:
	if ((fsm_stall == 1'd0) && (main_while_cond_i_cmp_i == 1'd1))
		next_state = LEGUP_F_main_BB_mmc_exit_loopexit_6;
	else if ((fsm_stall == 1'd0) && (main_while_cond_i_cmp_i == 1'd0))
		next_state = LEGUP_F_main_BB_while_body_i_3;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if ((((cur_state == LEGUP_0) & (fsm_stall == 1'd0)) & (start == 1'd1))) begin
		main_while_body_lr_ph_i_indvar3 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_else_i_5) & (fsm_stall == 1'd0)) & (main_if_else_i_cmp10_i == 1'd0))) */ begin
		main_while_body_lr_ph_i_indvar3 = main_if_else_i_indvar_next4;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_0) & (fsm_stall == 1'd0)) & (start == 1'd1))) begin
		main_while_body_lr_ph_i_indvar3_reg <= main_while_body_lr_ph_i_indvar3;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_else_i_5) & (fsm_stall == 1'd0)) & (main_if_else_i_cmp10_i == 1'd0))) begin
		main_while_body_lr_ph_i_indvar3_reg <= main_while_body_lr_ph_i_indvar3;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_0) & (fsm_stall == 1'd0)) & (start == 1'd1))) begin
		main_while_body_lr_ph_i_F2_0_ph15_i = 32'd7;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_else_i_5) & (fsm_stall == 1'd0)) & (main_if_else_i_cmp10_i == 1'd0))) */ begin
		main_while_body_lr_ph_i_F2_0_ph15_i = main_while_body_i_F2_011_i_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_0) & (fsm_stall == 1'd0)) & (start == 1'd1))) begin
		main_while_body_lr_ph_i_F2_0_ph15_i_reg <= main_while_body_lr_ph_i_F2_0_ph15_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_else_i_5) & (fsm_stall == 1'd0)) & (main_if_else_i_cmp10_i == 1'd0))) begin
		main_while_body_lr_ph_i_F2_0_ph15_i_reg <= main_while_body_lr_ph_i_F2_0_ph15_i;
	end
end
always @(*) begin
		main_while_body_lr_ph_i_bit_select3 = main_while_body_lr_ph_i_indvar3_reg[30:0];
end
always @(*) begin
		main_while_body_lr_ph_i_bit_select1 = main_while_body_lr_ph_i_indvar3_reg[29:0];
end
always @(*) begin
		main_while_body_lr_ph_i_bit_concat4 = {main_while_body_lr_ph_i_bit_select3[30:0], main_while_body_lr_ph_i_bit_concat4_bit_select_operand_2};
end
always @(*) begin
		main_while_body_lr_ph_i_bit_concat2 = {main_while_body_lr_ph_i_bit_select1[29:0], main_while_body_lr_ph_i_bit_concat2_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_while_body_lr_ph_i_sr_add = (main_while_body_lr_ph_i_bit_concat4 + main_while_body_lr_ph_i_bit_concat2);
end
always @(*) begin
		main_while_body_lr_ph_i_add2_i = (main_while_body_lr_ph_i_sr_add + 32'd12);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_lr_ph_i_1)) begin
		main_while_body_lr_ph_i_add2_i_reg <= main_while_body_lr_ph_i_add2_i;
	end
end
always @(*) begin
		main_while_body_lr_ph_i_F1_0_ph14_i = (main_while_body_lr_ph_i_sr_add + 32'd6);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_lr_ph_i_1)) begin
		main_while_body_lr_ph_i_F1_0_ph14_i_reg <= main_while_body_lr_ph_i_F1_0_ph14_i;
	end
end
always @(*) begin
		main_while_body_lr_ph_i_0 = (main_while_body_lr_ph_i_F2_0_ph15_i_reg + 32'd7);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_lr_ph_i_1)) begin
		main_while_body_lr_ph_i_0_reg <= main_while_body_lr_ph_i_0;
	end
end
always @(*) begin
		main_while_cond_i_add_i = (main_while_body_lr_ph_i_0_reg + main_while_body_i_sr_add7_reg);
end
always @(*) begin
		main_while_cond_i_cmp_i = (main_while_body_lr_ph_i_F1_0_ph14_i_reg == main_while_cond_i_add_i);
end
always @(*) begin
		main_while_cond_i_indvar_next = (main_while_body_i_indvar_reg + 32'd1);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_lr_ph_i_1) & (fsm_stall == 1'd0))) begin
		main_while_body_i_indvar = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_while_cond_i_2) & (fsm_stall == 1'd0)) & (main_while_cond_i_cmp_i == 1'd0))) */ begin
		main_while_body_i_indvar = main_while_cond_i_indvar_next;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_lr_ph_i_1) & (fsm_stall == 1'd0))) begin
		main_while_body_i_indvar_reg <= main_while_body_i_indvar;
	end
	if ((((cur_state == LEGUP_F_main_BB_while_cond_i_2) & (fsm_stall == 1'd0)) & (main_while_cond_i_cmp_i == 1'd0))) begin
		main_while_body_i_indvar_reg <= main_while_body_i_indvar;
	end
end
always @(*) begin
		main_while_body_i_bit_select = main_while_body_i_indvar_reg[28:0];
end
always @(*) begin
		main_while_body_i_sr_negate = (32'd0 - main_while_body_i_indvar_reg);
end
always @(*) begin
		main_while_body_i_bit_concat = {main_while_body_i_bit_select[28:0], main_while_body_i_bit_concat_bit_select_operand_2[2:0]};
end
always @(*) begin
		main_while_body_i_sr_add7 = (main_while_body_i_sr_negate + main_while_body_i_bit_concat);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i_3)) begin
		main_while_body_i_sr_add7_reg <= main_while_body_i_sr_add7;
	end
end
always @(*) begin
		main_while_body_i_F2_011_i = (main_while_body_lr_ph_i_F2_0_ph15_i_reg + main_while_body_i_sr_add7);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i_3)) begin
		main_while_body_i_F2_011_i_reg <= main_while_body_i_F2_011_i;
	end
end
always @(*) begin
		main_while_body_i_cmp1_i = ($signed(main_while_body_lr_ph_i_F1_0_ph14_i_reg) > $signed(main_while_body_i_F2_011_i_reg));
end
always @(*) begin
		main_if_else_i_cmp10_i = (main_while_body_lr_ph_i_add2_i_reg == main_while_body_i_F2_011_i_reg);
end
always @(*) begin
		main_if_else_i_indvar_next4 = (main_while_body_lr_ph_i_indvar3_reg + 32'd1);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_mmc_exit_loopexit_6) & (fsm_stall == 1'd0))) begin
		main_mmc_exit_F1_0_ph_lcssa_i = main_while_body_lr_ph_i_F1_0_ph14_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_mmc_exit_loopexit1_7) & (fsm_stall == 1'd0))) */ begin
		main_mmc_exit_F1_0_ph_lcssa_i = main_while_body_lr_ph_i_add2_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_mmc_exit_loopexit_6) & (fsm_stall == 1'd0))) begin
		main_mmc_exit_F1_0_ph_lcssa_i_reg <= main_mmc_exit_F1_0_ph_lcssa_i;
	end
	if (((cur_state == LEGUP_F_main_BB_mmc_exit_loopexit1_7) & (fsm_stall == 1'd0))) begin
		main_mmc_exit_F1_0_ph_lcssa_i_reg <= main_mmc_exit_F1_0_ph_lcssa_i;
	end
end
assign main_while_body_lr_ph_i_bit_concat4_bit_select_operand_2 = 1'd0;
assign main_while_body_lr_ph_i_bit_concat2_bit_select_operand_2 = 2'd0;
assign main_while_body_i_bit_concat_bit_select_operand_2 = 3'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_mmc_exit_8)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_mmc_exit_8)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "CycloneIV",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
