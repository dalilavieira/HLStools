library verilog;
use verilog.vl_types.all;
entity main is
    generic(
        LEGUP_0         : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LEGUP_F_main_BB_bb3_3_1: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        LEGUP_F_main_BB_bb3_3_2: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        LEGUP_F_main_BB_bb3_3_3: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        LEGUP_F_main_BB_bb3_3_4: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        LEGUP_F_main_BB_bb3_3_5: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        LEGUP_F_main_BB_bb3_3_7: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        LEGUP_F_main_BB_bb3_3_9: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        LEGUP_F_main_BB_bb3_3_11: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        LEGUP_F_main_BB_bb3_3_13: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        LEGUP_F_main_BB_bb3_3_14: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        LEGUP_F_main_BB_bb3_3_15: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        LEGUP_F_main_BB_bb3_3_17: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        LEGUP_F_main_BB_bb3_3_18: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        LEGUP_F_main_BB_bb3_3_19: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        LEGUP_F_main_BB_bb3_3_21: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        LEGUP_F_main_BB_bb3_3_22: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        LEGUP_F_main_BB_bb3_3_23: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        LEGUP_F_main_BB_bb3_3_25: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        LEGUP_F_main_BB_bb3_3_26: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        LEGUP_F_main_BB_bb3_3_27: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        LEGUP_F_main_BB_bb3_3_29: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        LEGUP_F_main_BB_bb15_30: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        LEGUP_F_main_BB_bb16_31: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        LEGUP_F_main_BB_return_32: vl_logic_vector(5 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        LEGUP_function_call_6: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        LEGUP_function_call_8: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        LEGUP_function_call_10: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        LEGUP_function_call_12: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        LEGUP_function_call_16: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        LEGUP_function_call_20: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        LEGUP_function_call_24: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        LEGUP_function_call_28: vl_logic_vector(5 downto 0) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0)
    );
    port(
        clk             : in     vl_logic;
        clk2x           : in     vl_logic;
        clk1x_follower  : in     vl_logic;
        reset           : in     vl_logic;
        start           : in     vl_logic;
        finish          : out    vl_logic;
        return_val      : out    vl_logic_vector(31 downto 0);
        memory_controller_enable_arbiter_a: out    vl_logic;
        memory_controller_address_arbiter_a: out    vl_logic_vector(31 downto 0);
        memory_controller_write_enable_arbiter_a: out    vl_logic;
        memory_controller_in_arbiter_a: out    vl_logic_vector(63 downto 0);
        memory_controller_size_arbiter_a: out    vl_logic_vector(1 downto 0);
        memory_controller_out_arbiter_a: in     vl_logic_vector(63 downto 0);
        memory_controller_enable_arbiter_b: out    vl_logic;
        memory_controller_address_arbiter_b: out    vl_logic_vector(31 downto 0);
        memory_controller_write_enable_arbiter_b: out    vl_logic;
        memory_controller_in_arbiter_b: out    vl_logic_vector(63 downto 0);
        memory_controller_size_arbiter_b: out    vl_logic_vector(1 downto 0);
        memory_controller_out_arbiter_b: in     vl_logic_vector(63 downto 0);
        memory_controller_waitrequest_arbiter: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LEGUP_0 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_1 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_2 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_3 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_4 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_5 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_7 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_9 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_11 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_13 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_14 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_15 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_17 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_18 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_19 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_21 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_22 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_23 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_25 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_26 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_27 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb3_3_29 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb15_30 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_bb16_31 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_F_main_BB_return_32 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_6 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_8 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_10 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_12 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_16 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_20 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_24 : constant is 2;
    attribute mti_svvh_generic_type of LEGUP_function_call_28 : constant is 2;
end main;
